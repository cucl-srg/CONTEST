***  Written by Yury Audzevich
*** 
***  Comments, suggestions for improvement and criticism welcome
***  E-mail:  yury.audzevich~at~cl.cam.ac.uk
*** 
*** 
***  Copyright 2003-2013, University of Cambridge, Computer Laboratory. 
***  Copyright and related rights are licensed under the Hardware License, 
***  Version 2.0 (the "License"); you may not use this file except in 
***  compliance with the License. You may obtain a copy of the License at
***  http://www.cl.cam.ac.uk/research/srg/netos/greenict/projects/contest/. 
***  Unless required by applicable law or agreed to in writing, software, 
***  hardware and materials distributed under this License is distributed 
***  on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
***  either express or implied. See the License for the specific language
***  governing permissions and limitations under the License.
*** 
*** 


***** HSPICE simulation using standard cell library  transistors *****
*** Noise margin for MCML gates ***

***** 45nm predictive technology model (FreePDK v1.4),  Typical conditions, 1.1V, 25C *****
.include "cells.spi"
.include "params.spi"

**** ================================================= ***
*** OPTIONS ***
.option post
.option nomod
.option co=255
*.option brief
.option dcon=1
.option lis_new=1
**.option captab 
.option accurate


**** ================================================= ***
*** MCML PARAMETERS ***
*** limits on the rotated curve
.param U = 0
.param UL = '-PARAM_MCML_SWING/sqrt(2)'
.param UH = 'PARAM_MCML_SWING/sqrt(2)'

************************************
*** Standard run without optimisation
.dc U UL UH 0.1m

************************************

**** ================================================= ***
*** MCML and ideal bias supplies
Vvdd VDD 0 PARAM_VDD_VOLTAGE
Vsss VSS 0 PARAM_VSS_VOLTAGE
*
Vvrefn VREFN 0 SWEEP_N_BIAS_VOLTAGE
Vvrefp VREFP 0 SWEEP_P_BIAS_VOLTAGE


*** For the methodology used please refer to the following source: 
*** F.J. List "The static noise margin of SRAM cells" 

**** ================================================= ***
*** Topology - single MCML INV instance
*** MCML INV requires Vin+ / Vin- signals generated simultaneously, 
*** so one instance of INV is sufficient for the analysis

Xinv1 Ip In Op On VDD VSS VREFP VREFN INV

*** Add small parasitic loads on outputs to be more realistic
C1 Op 0 CLOAD
C2 On 0 CLOAD

**** ================================================= ***
*** changing coordinates in 45 degree angle for Vin+ and Vin-
*** supply X = F(U,V)
EIp Ip VSS VOL = '(1/sqrt(2))*U + (1/sqrt(2))*V(V1p)'
EIn In VSS VOL = '-(1/sqrt(2))*U + (1/sqrt(2))*V(V1n)'

*** measure V = F(U,Y)
EV1p V1p VSS VOL = 'U + sqrt(2)*V(On)' 
EV1n V1n VSS VOL = '-U + sqrt(2)*V(Op)' 

*** create 2 complementary waveforms for '0->1' & '1->0' transitions
EV1d V1d 0 VOL = 'V(V1p) - V(V1n)'
EV2d V2d 0 VOL = 'V(V1n) - V(V1p)'

*** measure noise margin
EVD VD 0 VOL = 'ABS(V(V1d)-V(V2d))'

**** ================================================= ***
*** Measurements ***
**** ================================================= ***

*** Record the parameters in the .mt0 file
.meas DELIM0 param='0.0'
.meas dc result_vdd param='PARAM_VDD_VOLTAGE'
.meas dc result_vss param='PARAM_VSS_VOLTAGE'
.meas dc result_pulldown_width param='SWEEP_N_WIDTH'
.meas dc result_pulldown_length param='SWEEP_N_LENGTH'
.meas dc result_pullup_width param='SWEEP_P_WIDTH'
.meas dc result_pullup_length param='SWEEP_P_LENGTH'
.meas dc result_sink_width param='PARAM_NSOURCE_WIDTH'
.meas dc result_sink_length param='PARAM_NSOURCE_LENGTH'
.meas dc result_n_bias param='SWEEP_N_BIAS_VOLTAGE'
.meas dc result_p_bias param='SWEEP_P_BIAS_VOLTAGE'
.meas DELIM3 param='0.0'
.meas DELIM4 param='0.0'
.meas DELIM5 param='0.0'
.meas dc result_voltage_swing param='PARAM_MCML_SWING'
.meas dc MAXVD MAX V(VD)
.meas dc NOISE_MARGIN param='1/sqrt(2)*MAXVD'
.meas dc NM_PERCENT_OF_VSWING param='(NOISE_MARGIN/PARAM_MCML_SWING)*100'
