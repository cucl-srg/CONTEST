***  Written by Yury Audzevich
*** 
***  Comments, suggestions for improvement and criticism welcome
***  E-mail:  yury.audzevich~at~cl.cam.ac.uk
*** 
*** 
***  Copyright 2003-2013, University of Cambridge, Computer Laboratory. 
***  Copyright and related rights are licensed under the Hardware License, 
***  Version 2.0 (the "License"); you may not use this file except in 
***  compliance with the License. You may obtain a copy of the License at
***  http://www.cl.cam.ac.uk/research/srg/netos/greenict/projects/contest/. 
***  Unless required by applicable law or agreed to in writing, software, 
***  hardware and materials distributed under this License is distributed 
***  on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
***  either express or implied. See the License for the specific language
***  governing permissions and limitations under the License.
*** 
*** 


***** HSPICE simulation using standard cell library  transistors *****

***** 45nm predictive technology model (FreePDK v1.4),  Typical conditions, 1.1V, 25C *****
.include "/usr/groups/ecad/kits/commercial45_v2010_12/n45-hspice-model-TT_1V10_25.spi"

*********************************************************************
*** CMOS to MCML conversion circuit 
.subckt CMOS_to_MCML in outd outi mvdd vrfp vrfn cvdd gnda 
* CMOS INVs
M1 ini in gnda gnda NMOS_VTL W=SWEEP_CMOSN_WIDTH L=0.05U
M2 ini in cvdd cvdd PMOS_VTL W=SWEEP_CMOSP_WIDTH L=0.05U
*
M3 ind ini gnda gnda NMOS_VTL W=SWEEP_CMOSN_WIDTH L=0.05U
M4 ind ini cvdd cvdd PMOS_VTL W=SWEEP_CMOSP_WIDTH L=0.05U  
* MCML gate
M9 outi vrfp mvdd mvdd PMOS_VTL W=SWEEP_P_WIDTH L=SWEEP_P_LENGTH 
M10 outd vrfp mvdd mvdd PMOS_VTL W=SWEEP_P_WIDTH L=SWEEP_P_LENGTH 
M11 outi ind ic gnda NMOS_VTL W=SWEEP_N_WIDTH L=SWEEP_N_LENGTH
M12 outd ini ic gnda NMOS_VTL W=SWEEP_N_WIDTH L=SWEEP_N_LENGTH 
M13 ic vrfn gnda gnda NMOS_VTL W=PARAM_NSOURCE_WIDTH L=PARAM_NSOURCE_LENGTH
.ends CMOS_to_MCML


*********************************************************************
*** MCML to CMOS conversion
.subckt MCML_to_CMOS ind ini out mvdd vrfn gnda
* MCML gate
M1 mvdd pc pc mvdd PMOS_VTL W=SWEEP_P_WIDTH L=SWEEP_P_LENGTH
M2 mvdd nc nc mvdd PMOS_VTL W=SWEEP_P_WIDTH L=SWEEP_P_LENGTH
M3 ic ini pc gnda NMOS_VTL W=SWEEP_N_WIDTH L=SWEEP_N_LENGTH 
M4 ic ind nc gnda NMOS_VTL W=SWEEP_N_WIDTH L=SWEEP_N_LENGTH 
M5 gnda vrfn ic gnda NMOS_VTL W=PARAM_NSOURCE_WIDTH L=PARAM_NSOURCE_LENGTH
* CMOS INVs
M6 gnda bc bc gnda NMOS_VTL W=SWEEP_CMOSN_WIDTH L=0.05U
M7 mvdd nc bc mvdd PMOS_VTL W=SWEEP_CMOSP_WIDTH L=0.05U
*
M8 gnda bc ppa gnda NMOS_VTL W=SWEEP_CMOSN_WIDTH L=0.05U
M9 mvdd pc ppa mvdd PMOS_VTL W=SWEEP_CMOSP_WIDTH L=0.05U
*
M10 gnda ppa out gnda NMOS_VTL W=SWEEP_CMOSN_WIDTH L=0.05U
M11 mvdd ppa out mvdd PMOS_VTL W=SWEEP_CMOSP_WIDTH L=0.05U
.ends MCML_to_CMOS



*********************************************************************
*** MCML inverter - topological definition ***
.subckt INV An Ap Zn Zp VDD VSS VREFP VREFN
M1 Zn VREFP VDD VDD PMOS_VTL W=SWEEP_P_WIDTH L=SWEEP_P_LENGTH
M2 Zp VREFP VDD VDD PMOS_VTL W=SWEEP_P_WIDTH L=SWEEP_P_LENGTH
M3 Zn Ap nodeX VSS NMOS_VTL W=SWEEP_N_WIDTH L=SWEEP_N_LENGTH
M4 Zp An nodeX VSS NMOS_VTL W=SWEEP_N_WIDTH L=SWEEP_N_LENGTH
M5 nodeX VREFN VSS VSS NMOS_VTL W=PARAM_NSOURCE_WIDTH L=PARAM_NSOURCE_LENGTH
.ends INV



