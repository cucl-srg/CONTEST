***  Written by Yury Audzevich
*** 
***  Comments, suggestions for improvement and criticism welcome
***  E-mail:  yury.audzevich~at~cl.cam.ac.uk
*** 
*** 
***  Copyright 2003-2013, University of Cambridge, Computer Laboratory. 
***  Copyright and related rights are licensed under the Hardware License, 
***  Version 2.0 (the "License"); you may not use this file except in 
***  compliance with the License. You may obtain a copy of the License at
***  http://www.cl.cam.ac.uk/research/srg/netos/greenict/projects/contest/. 
***  Unless required by applicable law or agreed to in writing, software, 
***  hardware and materials distributed under this License is distributed 
***  on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
***  either express or implied. See the License for the specific language
***  governing permissions and limitations under the License.
*** 
*** 


*** 45nm predictive technology model (FreePDK v1.4),  Typical conditions, 1.1V, 25C ***

********************************************************************************
*** This file contains a collection of Design Parameters used in: 	     ***
*** optimization of douple-level MCML logic 				     ***	
********************************************************************************

*** MAIN PARAMETERS ***


*** Optimization ON/OFF ('1'/'0')  ***
.param OPT_PARAM_ON = 0

*** Gate under test (1) D-latch; (2) DFF+inv; (3) DFF-inv; (4) SEL;
*** (5) AND; (6) OR; (7) Other;
.param GATE_UND_TEST = 2

*** simulation time
.param PARAM_TIME_S = 0.1ps
.param PARAM_TIME_E = 6ns

*** measurement time
.param PARAM_MEAS_S = 100ps
.param PARAM_MEAS_E = 6ns

*** voltage swing ***
.param PARAM_MCML_SWING = 0.4
*.param PARAM_MCML_SWING = optw(0.2, 0.2, 0.45, 0.01)

*** level shifting ***
.param PARAM_MCML_LS = 'PARAM_MCML_SWING-(0.3*PARAM_MCML_SWING)'

*** supply voltages ***
.param PARAM_MCML_VDD_VOLTAGE = 0.9
.param PARAM_MCML_VSS_VOLTAGE = 0.0

*** derived parameters
.param PARAM_MCML_MID = '(PARAM_MCML_VDD_VOLTAGE + (PARAM_MCML_VDD_VOLTAGE-PARAM_MCML_SWING))/2'
.param PARAM_MCML_HALF_SWING = 'PARAM_MCML_SWING/2' 
.param PARAM_MCML_MIN = 'PARAM_MCML_VDD_VOLTAGE-PARAM_MCML_SWING'

*** parasitic capacitance
.param CLOAD = 0.05fF 

*** check for FANOUT ***
.param FANOUT_ON = 0

*** Define parameters to optimise and the ones to have fixed - the format is optw(initial, min, max, step)
*** In general HSPICE is more successful with fewer parameters to optimise when circuit has nonlinear responses to small deltas

*** Please comment/uncomment parameters that are needed for opt (2-4 parameters at a time for speed) ***
*** pull-up network
*.param SWEEP_P_WIDTH = optw(0.2U, 0.2U, 0.5U, 0.001U)
.param SWEEP_P_WIDTH=0.47U

*.param SWEEP_P_LENGTH = optw(0.1U, 0.1U, 0.15U, 0.005U)
.param SWEEP_P_LENGTH=0.11U

*** pull-down network
*.param SWEEP_N_WIDTH = optw(0.2U, 0.2U, 0.5U, 0.001U)
.param SWEEP_N_WIDTH=0.29U

*.param SWEEP_N_LENGTH = optw(lmin, lmin, 0.15U, 0.005U)
.param SWEEP_N_LENGTH= 0.05U

*** current sink 
.param PARAM_NSOURCE_WIDTH = 1.26U
*.param PARAM_NSOURCE_WIDTH = optw(1.0U, 1.0U, 3.0U, 0.001U)
*
.param PARAM_NSOURCE_LENGTH = 0.17U
*.param PARAM_NSOURCE_LENGTH = optw(lmin, lmin, 0.5U, 0.005U) 

*** level shifting current sink
.param PARAM_LS_N_WIDTH = 0.3U
*.param PARAM_LS_N_WIDTH = optw(0.2U, 0.2U, 5.0U, 0.001U)

.param PARAM_LS_N_LENGTH = 0.05U
*.param PARAM_LS_N_LENGTH = optw(lmin, lmin, 0.5U, 0.005U)

.param PARAM_LS_NS_WIDTH = 1.0U
*.param PARAM_LS_NS_WIDTH = optw(0.2U, 0.2U, 5.0U, 0.001U)

.param PARAM_LS_NS_LENGTH = 0.1U
*.param PARAM_LS_NS_LENGTH = optw(lmin, lmin, 0.5U, 0.005U) 
 

*** reference voltages
*.param SWEEP_N_BIAS_VOLTAGE = optw(0.3, 0.3, 0.7, 0.001)
.param SWEEP_N_BIAS_VOLTAGE = 0.55V

*.param SWEEP_P_BIAS_VOLTAGE = optw(20m, 20m, 300m , 0.1m)
.param SWEEP_P_BIAS_VOLTAGE = 50mV

*.param SWEEP_LEVEL_SHIFT_VOLTAGE = optw(0.01, 0.01, 0.35 , 0.001)
.param SWEEP_LEVEL_SHIFT_VOLTAGE = 0.1V

**** MAIN MCML INV params for testing ****
.param PARAM_INV_PW = 0.32U
.param PARAM_INV_PL = 0.07U

.param PARAM_INV_NW = 0.3U
.param PARAM_INV_NL = 'lmin'

.param PARAM_INV_NSW = 1.2U
.param PARAM_INV_NSL = 0.12U

.param PARAM_INV_VRP = 2mV
.param PARAM_INV_VRN = 0.53V


