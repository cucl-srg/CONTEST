***  Written by Yury Audzevich
*** 
***  Comments, suggestions for improvement and criticism welcome
***  E-mail:  yury.audzevich~at~cl.cam.ac.uk
*** 
*** 
***  Copyright 2003-2013, University of Cambridge, Computer Laboratory. 
***  Copyright and related rights are licensed under the Hardware License, 
***  Version 2.0 (the "License"); you may not use this file except in 
***  compliance with the License. You may obtain a copy of the License at
***  http://www.cl.cam.ac.uk/research/srg/netos/greenict/projects/contest/. 
***  Unless required by applicable law or agreed to in writing, software, 
***  hardware and materials distributed under this License is distributed 
***  on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
***  either express or implied. See the License for the specific language
***  governing permissions and limitations under the License.
*** 
*** 


***** HSPICE simulation using standard cell library  transistors *****
*** Noise margin for CMOS gates - testing approach specified below ***
*** Reference -- F.J. List, "The static noise margin of SRAM cells".  

***** 45nm predictive technology model (FreePDK v1.4),  Typical conditions, 1.1V, 25C *****
.include "/usr/groups/ecad/kits/commercial45_v2010_12/n45-hspice-model-TT_1V10_25.spi"

**** ================================================= ***
*** CMOS inverter ***
.subckt CMOS_INV IN OUT VDD VSS 
M1 OUT IN  VDD VDD PMOS_VTL W=CMOS_P_WIDTH L=CMOS_P_LENGTH
M2 OUT IN VSS VSS NMOS_VTL W=CMOS_N_WIDTH L=CMOS_N_LENGTH
.ends CMOS_INV

**** ================================================= ***
*** OPTIONS ***
.option post
.option nomod
.option co=255
*.option brief
.option dcon=1
.option lis_new=1
**.option captab 
.option accurate

**** ================================================= ***

*** parasitic capacitance
.param CLOAD = '0.05fF' 

******* CMOS SPECIFIC PARAMS ***********
* VDD & VSS
.param PARAM_CMOS_VDD = '1.1'
.param PARAM_CMOS_VSS = '0.0'

*** complementary pair
* P-type W & L
.param CMOS_P_WIDTH = 0.6U
.param CMOS_P_LENGTH = 'lmin'
* N-type W & L
.param CMOS_N_WIDTH = 0.2U
.param CMOS_N_LENGTH = 'lmin'
*
* rotated coordinate system (U,V)
** limits on U param variation
.param U = 0
.param UL = '-PARAM_CMOS_VDD/sqrt(2)'
.param UH = 'PARAM_CMOS_VDD/sqrt(2)'


************************************
*** Standard DC run without optimisation
.dc U UL UH 0.01

************************************

**** ================================================= ***
*** CMOS bias supplies 
Vvdd VDD 0 PARAM_CMOS_VDD
Vsss VSS 0 PARAM_CMOS_VSS

**** ================================================= ***
***************** CMOS testbench ******************
*** inv instances
Xi1 I1 O1 VDD VSS CMOS_INV	
Xi2 I2 O2 VDD VSS CMOS_INV

C1 O1 0 CLOAD
C2 O2 0 CLOAD

*** changing coordinates in 45 degree angle 
*** X and Y will have dependency on U and V as follows

*****************************************************
*** original function
EI1 I1 VSS VOL = '(1/sqrt(2))*U + (1/sqrt(2))*V(V1)'
EI2 I2 VSS VOL = '-(1/sqrt(2))*U + (1/sqrt(2))*V(V2)'

*** original function
EV1 V1 VSS VOL = 'U + sqrt(2)*V(O1)' 
EV2 V2 VSS VOL = '-U + sqrt(2)*V(O2)'

**** ================================================= ***
*** Measurements 
**** ================================================= ***
*** Record the parameters in the .mt0 file
.meas DELIM0 param='0.0'

EVD VDELTA 0 VOL = 'ABS(V(V1)-V(V2))'
.meas DC MAXD MAX V(VDELTA)
.meas DC SNM param='1/sqrt(2)*MAXD'



