*** 
***  Copyright 2003-2013, University of Cambridge, Computer Laboratory. 
***  Copyright and related rights are licensed under the Hardware License, 
***  Version 2.0 (the "License"); you may not use this file except in 
***  compliance with the License. You may obtain a copy of the License at
***  http://www.cl.cam.ac.uk/research/srg/netos/greenict/projects/contest/. 
***  Unless required by applicable law or agreed to in writing, software, 
***  hardware and materials distributed under this License is distributed 
***  on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
***  either express or implied. See the License for the specific language
***  governing permissions and limitations under the License.
*** 
*** 

*** SPICE structural netlist of 'SIPO4_64' after Design Compiler synthesis, based on port order in '/usr/groups/ecad/kits/commercial45_v2010_12/n45-library-netlist-noparasitics.spi' ***

.SUBCKT SIPO4_64 VDD_SIPO4_64 VSS_SIPO4_64 CLK_IN RESET_IN SERIAL_IN[0] SERIAL_IN[1] SERIAL_IN[2] SERIAL_IN[3] DATA_USED_OUT PARALLEL_OUT[0] PARALLEL_OUT[1] PARALLEL_OUT[2] PARALLEL_OUT[3] PARALLEL_OUT[4] PARALLEL_OUT[5] PARALLEL_OUT[6] PARALLEL_OUT[7] PARALLEL_OUT[8] PARALLEL_OUT[9] PARALLEL_OUT[10] PARALLEL_OUT[11] PARALLEL_OUT[12] PARALLEL_OUT[13] PARALLEL_OUT[14] PARALLEL_OUT[15] PARALLEL_OUT[16] PARALLEL_OUT[17] PARALLEL_OUT[18] PARALLEL_OUT[19] PARALLEL_OUT[20] PARALLEL_OUT[21] PARALLEL_OUT[22] PARALLEL_OUT[23] PARALLEL_OUT[24] PARALLEL_OUT[25] PARALLEL_OUT[26] PARALLEL_OUT[27] PARALLEL_OUT[28] PARALLEL_OUT[29] PARALLEL_OUT[30] PARALLEL_OUT[31] PARALLEL_OUT[32] PARALLEL_OUT[33] PARALLEL_OUT[34] PARALLEL_OUT[35] PARALLEL_OUT[36] PARALLEL_OUT[37] PARALLEL_OUT[38] PARALLEL_OUT[39] PARALLEL_OUT[40] PARALLEL_OUT[41] PARALLEL_OUT[42] PARALLEL_OUT[43] PARALLEL_OUT[44] PARALLEL_OUT[45] PARALLEL_OUT[46] PARALLEL_OUT[47] PARALLEL_OUT[48] PARALLEL_OUT[49] PARALLEL_OUT[50] PARALLEL_OUT[51] PARALLEL_OUT[52] PARALLEL_OUT[53] PARALLEL_OUT[54] PARALLEL_OUT[55] PARALLEL_OUT[56] PARALLEL_OUT[57] PARALLEL_OUT[58] PARALLEL_OUT[59] PARALLEL_OUT[60] PARALLEL_OUT[61] PARALLEL_OUT[62] PARALLEL_OUT[63]
*** instances
xpisos_0__SP1_16_shift_reg_reg_15_  SERIAL_IN[0]___rc n575___rc n585___rc pisos_0__SP1_16_shift_reg_15_ n91 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_14_  pisos_0__SP1_16_shift_reg_15____rc n577___rc n585___rc pisos_0__SP1_16_shift_reg_14_ n90 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_13_  pisos_0__SP1_16_shift_reg_14____rc n575___rc n585___rc pisos_0__SP1_16_shift_reg_13_ n89 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_12_  pisos_0__SP1_16_shift_reg_13____rc n575___rc n585___rc pisos_0__SP1_16_shift_reg_12_ n88 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_11_  pisos_0__SP1_16_shift_reg_12____rc n575___rc n585___rc pisos_0__SP1_16_shift_reg_11_ n87 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_10_  pisos_0__SP1_16_shift_reg_11____rc n575___rc n585___rc pisos_0__SP1_16_shift_reg_10_ n86 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_9_  pisos_0__SP1_16_shift_reg_10____rc n575___rc n585___rc pisos_0__SP1_16_shift_reg_9_ n85 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_8_  pisos_0__SP1_16_shift_reg_9____rc n576___rc n585___rc pisos_0__SP1_16_shift_reg_8_ n84 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_7_  pisos_0__SP1_16_shift_reg_8____rc n575___rc n585___rc pisos_0__SP1_16_shift_reg_7_ n83 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_6_  pisos_0__SP1_16_shift_reg_7____rc n577___rc n585___rc pisos_0__SP1_16_shift_reg_6_ n82 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_5_  pisos_0__SP1_16_shift_reg_6____rc n577___rc n585___rc pisos_0__SP1_16_shift_reg_5_ n81 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_4_  pisos_0__SP1_16_shift_reg_5____rc n577___rc n585___rc pisos_0__SP1_16_shift_reg_4_ n80 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_3_  pisos_0__SP1_16_shift_reg_4____rc n577___rc n585___rc pisos_0__SP1_16_shift_reg_3_ n79 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_2_  pisos_0__SP1_16_shift_reg_3____rc n577___rc n585___rc pisos_0__SP1_16_shift_reg_2_ n78 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_1_  pisos_0__SP1_16_shift_reg_2____rc n577___rc n585___rc pisos_0__SP1_16_shift_reg_1_ n77 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_shift_reg_reg_0_  pisos_0__SP1_16_shift_reg_1____rc n575___rc n585___rc SPICE_NETLIST_UNCONNECTED_1 n74 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_15_  SERIAL_IN[1]___rc n576___rc n585___rc pisos_1__SP1_16_shift_reg_15_ n109 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_14_  pisos_1__SP1_16_shift_reg_15____rc n577___rc n585___rc pisos_1__SP1_16_shift_reg_14_ n108 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_13_  pisos_1__SP1_16_shift_reg_14____rc n576___rc n585___rc pisos_1__SP1_16_shift_reg_13_ n107 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_12_  pisos_1__SP1_16_shift_reg_13____rc n576___rc n585___rc pisos_1__SP1_16_shift_reg_12_ n106 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_11_  pisos_1__SP1_16_shift_reg_12____rc n576___rc n585___rc pisos_1__SP1_16_shift_reg_11_ n105 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_10_  pisos_1__SP1_16_shift_reg_11____rc n576___rc n585___rc pisos_1__SP1_16_shift_reg_10_ n104 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_9_  pisos_1__SP1_16_shift_reg_10____rc n577___rc n585___rc pisos_1__SP1_16_shift_reg_9_ n103 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_8_  pisos_1__SP1_16_shift_reg_9____rc n577___rc n585___rc pisos_1__SP1_16_shift_reg_8_ n102 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_7_  pisos_1__SP1_16_shift_reg_8____rc n576___rc n585___rc pisos_1__SP1_16_shift_reg_7_ n101 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_6_  pisos_1__SP1_16_shift_reg_7____rc n577___rc n585___rc pisos_1__SP1_16_shift_reg_6_ n100 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_5_  pisos_1__SP1_16_shift_reg_6____rc n576___rc n585___rc pisos_1__SP1_16_shift_reg_5_ n99 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_4_  pisos_1__SP1_16_shift_reg_5____rc n576___rc n585___rc pisos_1__SP1_16_shift_reg_4_ n98 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_3_  pisos_1__SP1_16_shift_reg_4____rc n575___rc n585___rc pisos_1__SP1_16_shift_reg_3_ n97 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_2_  pisos_1__SP1_16_shift_reg_3____rc n576___rc n585___rc pisos_1__SP1_16_shift_reg_2_ n96 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_1_  pisos_1__SP1_16_shift_reg_2____rc n577___rc n585___rc pisos_1__SP1_16_shift_reg_1_ n95 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_shift_reg_reg_0_  pisos_1__SP1_16_shift_reg_1____rc n575___rc n585___rc SPICE_NETLIST_UNCONNECTED_2 n92 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_15_  SERIAL_IN[2]___rc n576___rc n584___rc pisos_2__SP1_16_shift_reg_15_ n127 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_14_  pisos_2__SP1_16_shift_reg_15____rc n572___rc n584___rc pisos_2__SP1_16_shift_reg_14_ n126 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_13_  pisos_2__SP1_16_shift_reg_14____rc n573___rc n584___rc pisos_2__SP1_16_shift_reg_13_ n125 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_12_  pisos_2__SP1_16_shift_reg_13____rc n572___rc n584___rc pisos_2__SP1_16_shift_reg_12_ n124 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_11_  pisos_2__SP1_16_shift_reg_12____rc n572___rc n584___rc pisos_2__SP1_16_shift_reg_11_ n123 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_10_  pisos_2__SP1_16_shift_reg_11____rc n574___rc n584___rc pisos_2__SP1_16_shift_reg_10_ n122 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_9_  pisos_2__SP1_16_shift_reg_10____rc n574___rc n584___rc pisos_2__SP1_16_shift_reg_9_ n121 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_8_  pisos_2__SP1_16_shift_reg_9____rc n574___rc n584___rc pisos_2__SP1_16_shift_reg_8_ n120 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_7_  pisos_2__SP1_16_shift_reg_8____rc n574___rc n584___rc pisos_2__SP1_16_shift_reg_7_ n119 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_6_  pisos_2__SP1_16_shift_reg_7____rc n574___rc n584___rc pisos_2__SP1_16_shift_reg_6_ n118 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_5_  pisos_2__SP1_16_shift_reg_6____rc n572___rc n584___rc pisos_2__SP1_16_shift_reg_5_ n117 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_4_  pisos_2__SP1_16_shift_reg_5____rc n573___rc n584___rc pisos_2__SP1_16_shift_reg_4_ n116 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_3_  pisos_2__SP1_16_shift_reg_4____rc n574___rc n584___rc pisos_2__SP1_16_shift_reg_3_ n115 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_2_  pisos_2__SP1_16_shift_reg_3____rc n573___rc n584___rc pisos_2__SP1_16_shift_reg_2_ n114 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_1_  pisos_2__SP1_16_shift_reg_2____rc n575___rc n584___rc pisos_2__SP1_16_shift_reg_1_ n113 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_shift_reg_reg_0_  pisos_2__SP1_16_shift_reg_1____rc n569___rc n584___rc SPICE_NETLIST_UNCONNECTED_3 n110 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_ctr_reg_1_  pisos_0__SP1_16_N2___rc n569___rc n584___rc pisos_0__SP1_16_ctr_1_ SPICE_NETLIST_UNCONNECTED_4 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_ctr_reg_2_  pisos_0__SP1_16_N3___rc n569___rc n584___rc pisos_0__SP1_16_ctr_2_ SPICE_NETLIST_UNCONNECTED_5 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_ctr_reg_3_  pisos_0__SP1_16_N4___rc n572___rc n584___rc pisos_0__SP1_16_ctr_3_ SPICE_NETLIST_UNCONNECTED_6 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_0_  n209___rc n569___rc n584___rc PARALLEL_OUT[0] SPICE_NETLIST_UNCONNECTED_7 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_1_  n208___rc n569___rc n584___rc PARALLEL_OUT[4] SPICE_NETLIST_UNCONNECTED_8 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_2_  n207___rc n569___rc n584___rc PARALLEL_OUT[8] SPICE_NETLIST_UNCONNECTED_9 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_3_  n206___rc n569___rc n584___rc PARALLEL_OUT[12] SPICE_NETLIST_UNCONNECTED_10 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_4_  n205___rc n569___rc n584___rc PARALLEL_OUT[16] SPICE_NETLIST_UNCONNECTED_11 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_5_  n204___rc n572___rc n583___rc PARALLEL_OUT[20] SPICE_NETLIST_UNCONNECTED_12 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_6_  n203___rc n572___rc n583___rc PARALLEL_OUT[24] SPICE_NETLIST_UNCONNECTED_13 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_7_  n202___rc n572___rc n583___rc PARALLEL_OUT[28] SPICE_NETLIST_UNCONNECTED_14 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_8_  n201___rc n572___rc n583___rc PARALLEL_OUT[32] SPICE_NETLIST_UNCONNECTED_15 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_9_  n200___rc n572___rc n583___rc PARALLEL_OUT[36] SPICE_NETLIST_UNCONNECTED_16 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_10_  n199___rc n572___rc n583___rc PARALLEL_OUT[40] SPICE_NETLIST_UNCONNECTED_17 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_11_  n198___rc n572___rc n583___rc PARALLEL_OUT[44] SPICE_NETLIST_UNCONNECTED_18 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_12_  n197___rc n572___rc n583___rc PARALLEL_OUT[48] SPICE_NETLIST_UNCONNECTED_19 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_13_  n196___rc n573___rc n583___rc PARALLEL_OUT[52] SPICE_NETLIST_UNCONNECTED_20 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_14_  n195___rc n572___rc n583___rc PARALLEL_OUT[56] SPICE_NETLIST_UNCONNECTED_21 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_0__SP1_16_PARALLEL_OUT_reg_15_  n194___rc n572___rc n583___rc PARALLEL_OUT[60] SPICE_NETLIST_UNCONNECTED_22 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_ctr_reg_1_  pisos_1__SP1_16_N2___rc n573___rc n583___rc pisos_1__SP1_16_ctr_1_ SPICE_NETLIST_UNCONNECTED_23 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_ctr_reg_2_  pisos_1__SP1_16_N3___rc n572___rc n584___rc pisos_1__SP1_16_ctr_2_ SPICE_NETLIST_UNCONNECTED_24 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_ctr_reg_3_  pisos_1__SP1_16_N4___rc n573___rc n584___rc pisos_1__SP1_16_ctr_3_ SPICE_NETLIST_UNCONNECTED_25 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_0_  n193___rc n572___rc n584___rc PARALLEL_OUT[1] SPICE_NETLIST_UNCONNECTED_26 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_1_  n192___rc n574___rc n584___rc PARALLEL_OUT[5] SPICE_NETLIST_UNCONNECTED_27 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_2_  n191___rc n574___rc n584___rc PARALLEL_OUT[9] SPICE_NETLIST_UNCONNECTED_28 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_3_  n190___rc n574___rc n584___rc PARALLEL_OUT[13] SPICE_NETLIST_UNCONNECTED_29 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_4_  n189___rc n574___rc n584___rc PARALLEL_OUT[17] SPICE_NETLIST_UNCONNECTED_30 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_5_  n188___rc n574___rc n584___rc PARALLEL_OUT[21] SPICE_NETLIST_UNCONNECTED_31 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_6_  n187___rc n574___rc n584___rc PARALLEL_OUT[25] SPICE_NETLIST_UNCONNECTED_32 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_7_  n186___rc n574___rc n584___rc PARALLEL_OUT[29] SPICE_NETLIST_UNCONNECTED_33 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_8_  n185___rc n572___rc n584___rc PARALLEL_OUT[33] SPICE_NETLIST_UNCONNECTED_34 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_9_  n184___rc n574___rc n584___rc PARALLEL_OUT[37] SPICE_NETLIST_UNCONNECTED_35 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_10_  n183___rc n577___rc n583___rc PARALLEL_OUT[41] SPICE_NETLIST_UNCONNECTED_36 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_11_  n182___rc n573___rc n583___rc PARALLEL_OUT[45] SPICE_NETLIST_UNCONNECTED_37 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_12_  n181___rc n576___rc n583___rc PARALLEL_OUT[49] SPICE_NETLIST_UNCONNECTED_38 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_13_  n180___rc n573___rc n583___rc PARALLEL_OUT[53] SPICE_NETLIST_UNCONNECTED_39 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_14_  n179___rc n575___rc n583___rc PARALLEL_OUT[57] SPICE_NETLIST_UNCONNECTED_40 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_1__SP1_16_PARALLEL_OUT_reg_15_  n178___rc n573___rc n583___rc PARALLEL_OUT[61] SPICE_NETLIST_UNCONNECTED_41 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_ctr_reg_1_  pisos_2__SP1_16_N2___rc n576___rc n585___rc pisos_2__SP1_16_ctr_1_ SPICE_NETLIST_UNCONNECTED_42 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_ctr_reg_2_  pisos_2__SP1_16_N3___rc n576___rc n584___rc pisos_2__SP1_16_ctr_2_ SPICE_NETLIST_UNCONNECTED_43 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_ctr_reg_3_  pisos_2__SP1_16_N4___rc n575___rc n584___rc pisos_2__SP1_16_ctr_3_ SPICE_NETLIST_UNCONNECTED_44 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_0_  n177___rc n573___rc n583___rc PARALLEL_OUT[2] SPICE_NETLIST_UNCONNECTED_45 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_1_  n176___rc n573___rc n583___rc PARALLEL_OUT[6] SPICE_NETLIST_UNCONNECTED_46 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_2_  n175___rc n570___rc n583___rc PARALLEL_OUT[10] SPICE_NETLIST_UNCONNECTED_47 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_3_  n174___rc n572___rc n583___rc PARALLEL_OUT[14] SPICE_NETLIST_UNCONNECTED_48 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_4_  n173___rc n573___rc n583___rc PARALLEL_OUT[18] SPICE_NETLIST_UNCONNECTED_49 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_5_  n172___rc n572___rc n583___rc PARALLEL_OUT[22] SPICE_NETLIST_UNCONNECTED_50 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_6_  n171___rc n572___rc n583___rc PARALLEL_OUT[26] SPICE_NETLIST_UNCONNECTED_51 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_7_  n170___rc n572___rc n583___rc PARALLEL_OUT[30] SPICE_NETLIST_UNCONNECTED_52 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_8_  n169___rc n572___rc n583___rc PARALLEL_OUT[34] SPICE_NETLIST_UNCONNECTED_53 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_9_  n168___rc n573___rc n583___rc PARALLEL_OUT[38] SPICE_NETLIST_UNCONNECTED_54 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_10_  n167___rc n572___rc n583___rc PARALLEL_OUT[42] SPICE_NETLIST_UNCONNECTED_55 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_11_  n166___rc n572___rc n583___rc PARALLEL_OUT[46] SPICE_NETLIST_UNCONNECTED_56 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_12_  n165___rc n572___rc n583___rc PARALLEL_OUT[50] SPICE_NETLIST_UNCONNECTED_57 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_13_  n164___rc n573___rc n583___rc PARALLEL_OUT[54] SPICE_NETLIST_UNCONNECTED_58 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_14_  n163___rc n572___rc n583___rc PARALLEL_OUT[58] SPICE_NETLIST_UNCONNECTED_59 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_2__SP1_16_PARALLEL_OUT_reg_15_  n162___rc n570___rc n582___rc PARALLEL_OUT[62] SPICE_NETLIST_UNCONNECTED_60 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_ctr_reg_1_  pisos_3__SP1_16_N2___rc n577___rc n585___rc pisos_3__SP1_16_ctr_1_ SPICE_NETLIST_UNCONNECTED_61 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_ctr_reg_2_  pisos_3__SP1_16_N3___rc n576___rc n585___rc pisos_3__SP1_16_ctr_2_ SPICE_NETLIST_UNCONNECTED_62 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_ctr_reg_3_  pisos_3__SP1_16_N4___rc n575___rc n585___rc pisos_3__SP1_16_ctr_3_ SPICE_NETLIST_UNCONNECTED_63 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_15_  SERIAL_IN[3]___rc n570___rc n582___rc pisos_3__SP1_16_shift_reg_15_ n145 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_14_  pisos_3__SP1_16_shift_reg_15____rc n571___rc n582___rc pisos_3__SP1_16_shift_reg_14_ n144 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_13_  pisos_3__SP1_16_shift_reg_14____rc n571___rc n582___rc pisos_3__SP1_16_shift_reg_13_ n143 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_12_  pisos_3__SP1_16_shift_reg_13____rc n577___rc n585___rc pisos_3__SP1_16_shift_reg_12_ n142 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_11_  pisos_3__SP1_16_shift_reg_12____rc n576___rc n585___rc pisos_3__SP1_16_shift_reg_11_ n141 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_10_  pisos_3__SP1_16_shift_reg_11____rc n575___rc n582___rc pisos_3__SP1_16_shift_reg_10_ n140 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_9_  pisos_3__SP1_16_shift_reg_10____rc n577___rc n585___rc pisos_3__SP1_16_shift_reg_9_ n139 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_8_  pisos_3__SP1_16_shift_reg_9____rc n570___rc n582___rc pisos_3__SP1_16_shift_reg_8_ n138 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_7_  pisos_3__SP1_16_shift_reg_8____rc n571___rc n582___rc pisos_3__SP1_16_shift_reg_7_ n137 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_6_  pisos_3__SP1_16_shift_reg_7____rc n571___rc n582___rc pisos_3__SP1_16_shift_reg_6_ n136 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_5_  pisos_3__SP1_16_shift_reg_6____rc n571___rc n582___rc pisos_3__SP1_16_shift_reg_5_ n135 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_4_  pisos_3__SP1_16_shift_reg_5____rc n571___rc n582___rc pisos_3__SP1_16_shift_reg_4_ n134 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_3_  pisos_3__SP1_16_shift_reg_4____rc n571___rc n582___rc pisos_3__SP1_16_shift_reg_3_ n133 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_2_  pisos_3__SP1_16_shift_reg_3____rc n571___rc n582___rc pisos_3__SP1_16_shift_reg_2_ n132 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_1_  pisos_3__SP1_16_shift_reg_2____rc n571___rc n582___rc pisos_3__SP1_16_shift_reg_1_ n131 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_shift_reg_reg_0_  pisos_3__SP1_16_shift_reg_1____rc n571___rc n582___rc SPICE_NETLIST_UNCONNECTED_64 n128 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_0_  n161___rc n571___rc n582___rc PARALLEL_OUT[3] SPICE_NETLIST_UNCONNECTED_65 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_1_  n160___rc n571___rc n582___rc PARALLEL_OUT[7] SPICE_NETLIST_UNCONNECTED_66 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_2_  n159___rc n571___rc n582___rc PARALLEL_OUT[11] SPICE_NETLIST_UNCONNECTED_67 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_3_  n158___rc n571___rc n582___rc PARALLEL_OUT[15] SPICE_NETLIST_UNCONNECTED_68 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_4_  n157___rc n571___rc n582___rc PARALLEL_OUT[19] SPICE_NETLIST_UNCONNECTED_69 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_5_  n156___rc n570___rc n582___rc PARALLEL_OUT[23] SPICE_NETLIST_UNCONNECTED_70 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_6_  n155___rc n570___rc n582___rc PARALLEL_OUT[27] SPICE_NETLIST_UNCONNECTED_71 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_7_  n154___rc n570___rc n582___rc PARALLEL_OUT[31] SPICE_NETLIST_UNCONNECTED_72 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_8_  n153___rc n570___rc n582___rc PARALLEL_OUT[35] SPICE_NETLIST_UNCONNECTED_73 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_9_  n152___rc n570___rc n582___rc PARALLEL_OUT[39] SPICE_NETLIST_UNCONNECTED_74 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_10_  n151___rc n570___rc n582___rc PARALLEL_OUT[43] SPICE_NETLIST_UNCONNECTED_75 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_11_  n150___rc n570___rc n582___rc PARALLEL_OUT[47] SPICE_NETLIST_UNCONNECTED_76 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_12_  n149___rc n570___rc n582___rc PARALLEL_OUT[51] SPICE_NETLIST_UNCONNECTED_77 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_13_  n148___rc n570___rc n582___rc PARALLEL_OUT[55] SPICE_NETLIST_UNCONNECTED_78 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_14_  n147___rc n570___rc n582___rc PARALLEL_OUT[59] SPICE_NETLIST_UNCONNECTED_79 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xpisos_3__SP1_16_PARALLEL_OUT_reg_15_  n146___rc n570___rc n582___rc PARALLEL_OUT[63] SPICE_NETLIST_UNCONNECTED_80 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xU170  n231___rc n496___rc n322___rc n197 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU174  n562___rc n233___rc n234 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU243  n443___rc n354___rc pisos_1__SP1_16_N4 VDD_SIPO4_64 VSS_SIPO4_64  XNOR2_X1
xU244  pisos_1__SP1_16_ctr_2____rc n229___rc n284___rc n443 VDD_SIPO4_64 VSS_SIPO4_64  AND3_X1
xU245  n485___rc n284 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU298  n337___rc n492___rc n322 VDD_SIPO4_64 VSS_SIPO4_64  AND2_X4
xU305  n440___rc n328___rc pisos_0__SP1_16_N4 VDD_SIPO4_64 VSS_SIPO4_64  XNOR2_X1
xU306  n531___rc n328 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU307  n447___rc n492___rc n353___rc n440 VDD_SIPO4_64 VSS_SIPO4_64  NOR3_X1
xU309  n446___rc n361___rc pisos_2__SP1_16_N4 VDD_SIPO4_64 VSS_SIPO4_64  XNOR2_X1
xU311  n447___rc n468___rc n362___rc n446 VDD_SIPO4_64 VSS_SIPO4_64  NOR3_X1
xU312  n450___rc n363___rc pisos_3__SP1_16_N4 VDD_SIPO4_64 VSS_SIPO4_64  XNOR2_X1
xU314  n447___rc n451___rc n364___rc n450 VDD_SIPO4_64 VSS_SIPO4_64  NOR3_X1
xU333  n531___rc n352 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU334  pisos_1__SP1_16_ctr_3____rc n354 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU335  n349___rc pisos_1__SP1_16_ctr_1____rc n350 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU345  n529___rc n361 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU346  pisos_3__SP1_16_ctr_3____rc n363 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU369  n578___rc n135___rc n376 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU371  n578___rc n145___rc n367 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU373  n578___rc n131___rc n380 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU375  n578___rc n134___rc n377 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU377  n578___rc n141___rc n371 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU380  n578___rc n128___rc n381 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU382  n578___rc n138___rc n374 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU384  n578___rc n143___rc n369 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU386  n578___rc n133___rc n378 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU388  n578___rc n136___rc n375 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU390  n578___rc n140___rc n372 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU392  n578___rc n139___rc n373 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU394  n578___rc n142___rc n370 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU396  n578___rc n144___rc n368 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU397  n580___rc n117___rc n392 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU398  n580___rc n123___rc n387 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU399  n397___rc n489___rc n562___rc n183 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU400  n408___rc n503___rc n322___rc n204 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU401  n339___rc n81___rc n408 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU402  n580___rc n127___rc n383 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU403  n580___rc n126___rc n384 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU404  n406___rc n501___rc n322___rc n202 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU405  n339___rc n83___rc n406 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU406  n580___rc n114___rc n394 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU407  n580___rc n113___rc n395 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU408  n580___rc n118___rc n391 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU409  n410___rc n505___rc n322___rc n206 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU410  n339___rc n79___rc n410 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU411  n580___rc n110___rc n396 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU412  n580___rc n116___rc n393 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU413  n409___rc n504___rc n322___rc n205 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU414  n339___rc n80___rc n409 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU415  n580___rc n121___rc n389 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU416  n580___rc n122___rc n388 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU417  n413___rc n508___rc n322___rc n209 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU418  n339___rc n74___rc n413 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU419  n403___rc n498___rc n322___rc n199 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU420  n339___rc n86___rc n403 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU421  n407___rc n502___rc n322___rc n203 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU422  n339___rc n82___rc n407 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU423  n580___rc n124___rc n386 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU424  n580___rc n125___rc n385 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU425  n412___rc n507___rc n322___rc n208 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU426  n339___rc n77___rc n412 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU427  n402___rc n497___rc n322___rc n198 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU428  n339___rc n87___rc n402 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU429  n405___rc n500___rc n322___rc n201 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU430  n339___rc n84___rc n405 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU431  n399___rc n493___rc n322___rc n194 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU432  n339___rc n91___rc n399 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU433  n411___rc n506___rc n322___rc n207 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU434  n339___rc n78___rc n411 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU435  n580___rc n119___rc n390 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU436  n404___rc n499___rc n322___rc n200 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU437  n339___rc n85___rc n404 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU438  n400___rc n494___rc n322___rc n195 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU439  n401___rc n495___rc n322___rc n196 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU440  n339___rc n89___rc n401 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU441  pisos_3__SP1_16_ctr_0____rc n366___rc n365___rc DATA_USED_OUT VDD_SIPO4_64 VSS_SIPO4_64  AOI21_X1
xU454  n229___rc pisos_0__SP1_16_ctr_1____rc n492___rc n447___rc pisos_0__SP1_16_N2 VDD_SIPO4_64 VSS_SIPO4_64  AOI22_X1
xU456  n229___rc pisos_0__SP1_16_ctr_1____rc n438 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU457  n440___rc n353___rc n438___rc pisos_0__SP1_16_N3 VDD_SIPO4_64 VSS_SIPO4_64  AOI21_X1
xU458  n229___rc pisos_1__SP1_16_ctr_1____rc n485___rc n447___rc pisos_1__SP1_16_N2 VDD_SIPO4_64 VSS_SIPO4_64  AOI22_X1
xU460  n229___rc pisos_1__SP1_16_ctr_1____rc n441 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU461  n443___rc n355___rc n441___rc pisos_1__SP1_16_N3 VDD_SIPO4_64 VSS_SIPO4_64  AOI21_X1
xU462  n229___rc pisos_2__SP1_16_ctr_1____rc n468___rc n447___rc pisos_2__SP1_16_N2 VDD_SIPO4_64 VSS_SIPO4_64  AOI22_X1
xU464  n229___rc pisos_2__SP1_16_ctr_1____rc n444 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU465  n446___rc n362___rc n444___rc pisos_2__SP1_16_N3 VDD_SIPO4_64 VSS_SIPO4_64  AOI21_X1
xU466  n229___rc pisos_3__SP1_16_ctr_1____rc n451___rc n447___rc pisos_3__SP1_16_N2 VDD_SIPO4_64 VSS_SIPO4_64  AOI22_X1
xU468  n229___rc pisos_3__SP1_16_ctr_1____rc n448 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU469  n450___rc n364___rc n448___rc pisos_3__SP1_16_N3 VDD_SIPO4_64 VSS_SIPO4_64  AOI21_X1
xU502  PARALLEL_OUT[57]___rc n486 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU503  PARALLEL_OUT[53]___rc n487 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU504  PARALLEL_OUT[45]___rc n488 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU505  PARALLEL_OUT[41]___rc n489 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU506  PARALLEL_OUT[21]___rc n490 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU507  PARALLEL_OUT[5]___rc n491 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU508  PARALLEL_OUT[60]___rc n493 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU509  PARALLEL_OUT[56]___rc n494 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU510  PARALLEL_OUT[52]___rc n495 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU511  PARALLEL_OUT[48]___rc n496 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU512  PARALLEL_OUT[44]___rc n497 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU513  PARALLEL_OUT[40]___rc n498 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU514  PARALLEL_OUT[36]___rc n499 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU515  PARALLEL_OUT[32]___rc n500 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU516  PARALLEL_OUT[28]___rc n501 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU517  PARALLEL_OUT[24]___rc n502 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU518  PARALLEL_OUT[20]___rc n503 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU519  PARALLEL_OUT[16]___rc n504 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU520  PARALLEL_OUT[12]___rc n505 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU521  PARALLEL_OUT[8]___rc n506 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU522  PARALLEL_OUT[4]___rc n507 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU523  PARALLEL_OUT[0]___rc n508 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU212  n266___rc n264___rc n193 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU238  n283___rc n282___rc n192 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU217  n270___rc n268___rc n191 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU172  n234___rc n232___rc n190 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU182  n242___rc n240___rc n189 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU226  n274___rc n273___rc n188 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU192  n250___rc n248___rc n187 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU197  n254___rc n252___rc n186 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU187  n246___rc n244___rc n185 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU202  n258___rc n256___rc n184 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU232  n279___rc n278___rc n182 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU177  n238___rc n236___rc n181 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU229  n277___rc n276___rc n180 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU207  n262___rc n260___rc n178 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU275  n396___rc n305___rc n177 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU269  n395___rc n301___rc n176 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU266  n394___rc n299___rc n175 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU254  n290___rc n115___rc n580___rc n174 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU278  n393___rc n307___rc n173 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU250  n392___rc n288___rc n172 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU272  n391___rc n303___rc n171 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU293  n390___rc n317___rc n170 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU297  n319___rc n120___rc n580___rc n169 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU281  n389___rc n309___rc n168 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU284  n388___rc n311___rc n167 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU257  n387___rc n293___rc n166 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU287  n386___rc n313___rc n165 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU290  n385___rc n315___rc n164 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU263  n384___rc n297___rc n163 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU260  n383___rc n295___rc n162 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU171  n322___rc n358___rc n231 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU322  n322___rc n338___rc n400 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU216  n562___rc n265___rc n266 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU213  n562___rc n267___rc n264 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU236  n562___rc n323___rc n283 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU237  n491___rc n562___rc n282 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU221  n562___rc n269___rc n270 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU218  n562___rc n271___rc n268 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU173  n562___rc n235___rc n232 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU186  n562___rc n241___rc n242 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU183  n562___rc n243___rc n240 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU224  n562___rc n324___rc n274 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU225  n490___rc n562___rc n273 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU196  n562___rc n249___rc n250 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU193  n562___rc n251___rc n248 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU201  n562___rc n253___rc n254 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU198  n562___rc n255___rc n252 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU191  n562___rc n245___rc n246 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU188  n562___rc n247___rc n244 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU206  n562___rc n257___rc n258 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU203  n562___rc n259___rc n256 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU320  n562___rc n336___rc n397 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU230  n562___rc n326___rc n279 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU231  n488___rc n562___rc n278 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU181  n562___rc n237___rc n238 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU178  n562___rc n239___rc n236 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU227  n562___rc n327___rc n277 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU228  n487___rc n562___rc n276 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU233  n562___rc n325___rc n281 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU211  n562___rc n261___rc n262 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU208  n562___rc n263___rc n260 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU274  n580___rc PARALLEL_OUT[2]___rc n305 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU268  n580___rc PARALLEL_OUT[6]___rc n301 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU265  n580___rc PARALLEL_OUT[10]___rc n299 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU253  n580___rc PARALLEL_OUT[14]___rc n290 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU277  n580___rc PARALLEL_OUT[18]___rc n307 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU249  n580___rc PARALLEL_OUT[22]___rc n288 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU271  n580___rc PARALLEL_OUT[26]___rc n303 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU292  n580___rc PARALLEL_OUT[30]___rc n317 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU296  n580___rc PARALLEL_OUT[34]___rc n319 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU280  n580___rc PARALLEL_OUT[38]___rc n309 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU283  n580___rc PARALLEL_OUT[42]___rc n311 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU256  n580___rc PARALLEL_OUT[46]___rc n293 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU286  n580___rc PARALLEL_OUT[50]___rc n313 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU289  n580___rc PARALLEL_OUT[54]___rc n315 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU262  n580___rc PARALLEL_OUT[58]___rc n297 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU259  n580___rc PARALLEL_OUT[62]___rc n295 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU347  pisos_2__SP1_16_ctr_2____rc pisos_2__SP1_16_ctr_3____rc n359 VDD_SIPO4_64 VSS_SIPO4_64  NOR2_X1
xU344  n88___rc n358 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU321  n90___rc n338 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU215  n92___rc n265 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU214  PARALLEL_OUT[1]___rc n267 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU299  n95___rc n323 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU220  n96___rc n269 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU219  PARALLEL_OUT[9]___rc n271 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU176  n97___rc n233 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU175  PARALLEL_OUT[13]___rc n235 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU185  n98___rc n241 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU184  PARALLEL_OUT[17]___rc n243 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU300  n99___rc n324 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU195  n100___rc n249 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU194  PARALLEL_OUT[25]___rc n251 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU200  n101___rc n253 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU199  PARALLEL_OUT[29]___rc n255 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU190  n102___rc n245 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU189  PARALLEL_OUT[33]___rc n247 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU205  n103___rc n257 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU204  PARALLEL_OUT[37]___rc n259 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU319  n104___rc n336 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU302  n105___rc n326 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU180  n106___rc n237 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU179  PARALLEL_OUT[49]___rc n239 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU303  n107___rc n327 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU301  n108___rc n325 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU210  n109___rc n261 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU209  PARALLEL_OUT[61]___rc n263 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU242  pisos_3__SP1_16_ctr_0____rc n447 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU337  n348___rc pisos_0__SP1_16_ctr_1____rc n351 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU366  pisos_0__SP1_16_ctr_1____rc n492 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU336  pisos_0__SP1_16_ctr_2____rc pisos_0__SP1_16_ctr_3____rc n348 VDD_SIPO4_64 VSS_SIPO4_64  NOR2_X1
xU367  pisos_1__SP1_16_ctr_1____rc n485 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU350  pisos_2__SP1_16_ctr_2____rc n362 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU349  pisos_3__SP1_16_ctr_2____rc n364 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU341  pisos_0__SP1_16_ctr_2____rc n353 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU365  pisos_2__SP1_16_ctr_1____rc n468 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU364  pisos_3__SP1_16_ctr_1____rc n451 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU340  pisos_1__SP1_16_ctr_2____rc n355 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xpisos_3__SP1_16_ctr_reg_0_  pisos_3__SP1_16_N1___rc n569___rc n584___rc pisos_3__SP1_16_ctr_0_ pisos_3__SP1_16_N1 VDD_SIPO4_64 VSS_SIPO4_64  DFFR_X1
xU328  pisos_3__SP1_16_ctr_1____rc n360___rc n359___rc pisos_2__SP1_16_ctr_1____rc n365 VDD_SIPO4_64 VSS_SIPO4_64  AOI22_X1
xU348  pisos_3__SP1_16_ctr_2____rc pisos_3__SP1_16_ctr_3____rc n360 VDD_SIPO4_64 VSS_SIPO4_64  NOR2_X1
xU528  n517___rc n132___rc n578___rc n159 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU529  n527___rc n137___rc n578___rc n154 VDD_SIPO4_64 VSS_SIPO4_64  OAI21_X1
xU534  n578___rc PARALLEL_OUT[23]___rc n512 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU535  n512___rc n376___rc n156 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU536  n578___rc PARALLEL_OUT[63]___rc n513 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU537  n513___rc n367___rc n146 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU538  n578___rc PARALLEL_OUT[7]___rc n514 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU539  n514___rc n380___rc n160 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU540  n578___rc PARALLEL_OUT[19]___rc n515 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU541  n515___rc n377___rc n157 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU542  n578___rc PARALLEL_OUT[47]___rc n516 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU543  n516___rc n371___rc n150 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU544  n578___rc PARALLEL_OUT[11]___rc n517 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU545  n578___rc PARALLEL_OUT[3]___rc n518 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU546  n518___rc n381___rc n161 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU547  n578___rc PARALLEL_OUT[35]___rc n519 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU548  n519___rc n374___rc n153 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU549  n578___rc PARALLEL_OUT[55]___rc n520 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU550  n520___rc n369___rc n148 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU551  n578___rc PARALLEL_OUT[15]___rc n521 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU552  n521___rc n378___rc n158 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU553  n578___rc PARALLEL_OUT[27]___rc n522 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU554  n522___rc n375___rc n155 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU555  n578___rc PARALLEL_OUT[43]___rc n523 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU556  n523___rc n372___rc n151 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU557  n578___rc PARALLEL_OUT[39]___rc n524 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU558  n524___rc n373___rc n152 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU559  n578___rc PARALLEL_OUT[51]___rc n525 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU560  n525___rc n370___rc n149 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU561  n578___rc PARALLEL_OUT[59]___rc n526 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU562  n526___rc n368___rc n147 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU563  n578___rc PARALLEL_OUT[31]___rc n527 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU565  pisos_2__SP1_16_ctr_3____rc n529 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X1
xU566  n530___rc n366 VDD_SIPO4_64 VSS_SIPO4_64  INV_X1
xU567  n351___rc n350___rc n530 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU582  n567___rc n572 VDD_SIPO4_64 VSS_SIPO4_64  INV_X4
xU574  n568___rc n575 VDD_SIPO4_64 VSS_SIPO4_64  INV_X2
xU572  n568___rc n577 VDD_SIPO4_64 VSS_SIPO4_64  INV_X2
xU573  n568___rc n576 VDD_SIPO4_64 VSS_SIPO4_64  INV_X2
xU235  n281___rc n280___rc n179 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU581  n567___rc n573 VDD_SIPO4_64 VSS_SIPO4_64  INV_X2
xU530  n581___rc n583 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X4
xU526  n581___rc n585 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X4
xU533  n581___rc n582 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X4
xU591  n566___rc n569 VDD_SIPO4_64 VSS_SIPO4_64  INV_X2
xU576  n566___rc n574 VDD_SIPO4_64 VSS_SIPO4_64  INV_X4
xU584  n566___rc n571 VDD_SIPO4_64 VSS_SIPO4_64  INV_X4
xU585  n566___rc n570 VDD_SIPO4_64 VSS_SIPO4_64  INV_X4
xU588  RESET_IN___rc n566 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X4
xU568  n579___rc n580 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X4
xU241  n357___rc pisos_3__SP1_16_ctr_0____rc n337 VDD_SIPO4_64 VSS_SIPO4_64  AND2_X2
xU564  pisos_0__SP1_16_ctr_3____rc n531 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X2
xU583  RESET_IN___rc n567 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X2
xU575  RESET_IN___rc n568 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X2
xU527  n581___rc n584 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X8
xU166  pisos_3__SP1_16_ctr_0____rc n229 VDD_SIPO4_64 VSS_SIPO4_64  BUF_X2
xU338  pisos_1__SP1_16_ctr_2____rc pisos_1__SP1_16_ctr_3____rc n349 VDD_SIPO4_64 VSS_SIPO4_64  NOR2_X1
xU329  n362___rc pisos_3__SP1_16_ctr_0____rc n344 VDD_SIPO4_64 VSS_SIPO4_64  AND2_X1
xU531  n468___rc n361___rc n509 VDD_SIPO4_64 VSS_SIPO4_64  AND2_X2
xU343  n352___rc n353___rc n357 VDD_SIPO4_64 VSS_SIPO4_64  AND2_X2
xU234  n486___rc n562___rc n280 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X1
xU240  n337___rc n492___rc n339 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X4
xU317  n344___rc n509___rc n579 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X2
xU594  n354___rc pisos_3__SP1_16_ctr_0____rc n561 VDD_SIPO4_64 VSS_SIPO4_64  AND2_X2
xU595  CLK_IN___rc n564 VDD_SIPO4_64 VSS_SIPO4_64  INV_X2
xU596  n559___rc n560___rc n578 VDD_SIPO4_64 VSS_SIPO4_64  OR2_X4
xU597  n451___rc n363___rc n560 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU598  n364___rc pisos_3__SP1_16_ctr_0____rc n559 VDD_SIPO4_64 VSS_SIPO4_64  NAND2_X1
xU599  n561___rc n355___rc n485___rc n562 VDD_SIPO4_64 VSS_SIPO4_64  AND3_X4
xU600  n564___rc n581 VDD_SIPO4_64 VSS_SIPO4_64  INV_X4
*** Estimated net resistances from Design Compiler
r1 CLK_IN CLK_IN___rc 4.0
r2 DATA_USED_OUT DATA_USED_OUT___rc 39.0
r3 PARALLEL_OUT[0] PARALLEL_OUT[0]___rc 61.0
r4 PARALLEL_OUT[10] PARALLEL_OUT[10]___rc 68.0
r5 PARALLEL_OUT[11] PARALLEL_OUT[11]___rc 40.0
r6 PARALLEL_OUT[12] PARALLEL_OUT[12]___rc 53.0
r7 PARALLEL_OUT[13] PARALLEL_OUT[13]___rc 18.0
r8 PARALLEL_OUT[14] PARALLEL_OUT[14]___rc 42.0
r9 PARALLEL_OUT[15] PARALLEL_OUT[15]___rc 44.0
r10 PARALLEL_OUT[16] PARALLEL_OUT[16]___rc 25.0
r11 PARALLEL_OUT[17] PARALLEL_OUT[17]___rc 21.0
r12 PARALLEL_OUT[18] PARALLEL_OUT[18]___rc 47.0
r13 PARALLEL_OUT[19] PARALLEL_OUT[19]___rc 71.0
r14 PARALLEL_OUT[1] PARALLEL_OUT[1]___rc 59.0
r15 PARALLEL_OUT[20] PARALLEL_OUT[20]___rc 38.0
r16 PARALLEL_OUT[21] PARALLEL_OUT[21]___rc 37.0
r17 PARALLEL_OUT[22] PARALLEL_OUT[22]___rc 34.0
r18 PARALLEL_OUT[23] PARALLEL_OUT[23]___rc 60.0
r19 PARALLEL_OUT[24] PARALLEL_OUT[24]___rc 47.0
r20 PARALLEL_OUT[25] PARALLEL_OUT[25]___rc 63.0
r21 PARALLEL_OUT[26] PARALLEL_OUT[26]___rc 55.0
r22 PARALLEL_OUT[27] PARALLEL_OUT[27]___rc 65.0
r23 PARALLEL_OUT[28] PARALLEL_OUT[28]___rc 49.0
r24 PARALLEL_OUT[29] PARALLEL_OUT[29]___rc 46.0
r25 PARALLEL_OUT[2] PARALLEL_OUT[2]___rc 69.0
r26 PARALLEL_OUT[30] PARALLEL_OUT[30]___rc 46.0
r27 PARALLEL_OUT[31] PARALLEL_OUT[31]___rc 36.0
r28 PARALLEL_OUT[32] PARALLEL_OUT[32]___rc 61.0
r29 PARALLEL_OUT[33] PARALLEL_OUT[33]___rc 39.0
r30 PARALLEL_OUT[34] PARALLEL_OUT[34]___rc 59.0
r31 PARALLEL_OUT[35] PARALLEL_OUT[35]___rc 71.0
r32 PARALLEL_OUT[36] PARALLEL_OUT[36]___rc 42.0
r33 PARALLEL_OUT[37] PARALLEL_OUT[37]___rc 28.0
r34 PARALLEL_OUT[38] PARALLEL_OUT[38]___rc 22.0
r35 PARALLEL_OUT[39] PARALLEL_OUT[39]___rc 61.0
r36 PARALLEL_OUT[3] PARALLEL_OUT[3]___rc 61.0
r37 PARALLEL_OUT[40] PARALLEL_OUT[40]___rc 48.0
r38 PARALLEL_OUT[41] PARALLEL_OUT[41]___rc 72.0
r39 PARALLEL_OUT[42] PARALLEL_OUT[42]___rc 32.0
r40 PARALLEL_OUT[43] PARALLEL_OUT[43]___rc 52.0
r41 PARALLEL_OUT[44] PARALLEL_OUT[44]___rc 20.0
r42 PARALLEL_OUT[45] PARALLEL_OUT[45]___rc 67.0
r43 PARALLEL_OUT[46] PARALLEL_OUT[46]___rc 40.0
r44 PARALLEL_OUT[47] PARALLEL_OUT[47]___rc 60.0
r45 PARALLEL_OUT[48] PARALLEL_OUT[48]___rc 69.0
r46 PARALLEL_OUT[49] PARALLEL_OUT[49]___rc 100.0
r47 PARALLEL_OUT[4] PARALLEL_OUT[4]___rc 44.0
r48 PARALLEL_OUT[50] PARALLEL_OUT[50]___rc 43.0
r49 PARALLEL_OUT[51] PARALLEL_OUT[51]___rc 81.0
r50 PARALLEL_OUT[52] PARALLEL_OUT[52]___rc 87.0
r51 PARALLEL_OUT[53] PARALLEL_OUT[53]___rc 64.0
r52 PARALLEL_OUT[54] PARALLEL_OUT[54]___rc 34.0
r53 PARALLEL_OUT[55] PARALLEL_OUT[55]___rc 51.0
r54 PARALLEL_OUT[56] PARALLEL_OUT[56]___rc 44.0
r55 PARALLEL_OUT[57] PARALLEL_OUT[57]___rc 67.0
r56 PARALLEL_OUT[58] PARALLEL_OUT[58]___rc 38.0
r57 PARALLEL_OUT[59] PARALLEL_OUT[59]___rc 55.0
r58 PARALLEL_OUT[5] PARALLEL_OUT[5]___rc 23.0
r59 PARALLEL_OUT[60] PARALLEL_OUT[60]___rc 58.0
r60 PARALLEL_OUT[61] PARALLEL_OUT[61]___rc 72.0
r61 PARALLEL_OUT[62] PARALLEL_OUT[62]___rc 91.0
r62 PARALLEL_OUT[63] PARALLEL_OUT[63]___rc 35.0
r63 PARALLEL_OUT[6] PARALLEL_OUT[6]___rc 75.0
r64 PARALLEL_OUT[7] PARALLEL_OUT[7]___rc 54.0
r65 PARALLEL_OUT[8] PARALLEL_OUT[8]___rc 51.0
r66 PARALLEL_OUT[9] PARALLEL_OUT[9]___rc 38.0
r67 RESET_IN RESET_IN___rc 206.0
r68 SERIAL_IN[0] SERIAL_IN[0]___rc 11.0
r69 SERIAL_IN[1] SERIAL_IN[1]___rc 9.0
r70 SERIAL_IN[2] SERIAL_IN[2]___rc 7.0
r71 SERIAL_IN[3] SERIAL_IN[3]___rc 44.0
r72 n100 n100___rc 98.0
r73 n101 n101___rc 55.0
r74 n102 n102___rc 29.0
r75 n103 n103___rc 36.0
r76 n104 n104___rc 26.0
r77 n105 n105___rc 14.0
r78 n106 n106___rc 82.0
r79 n107 n107___rc 38.0
r80 n108 n108___rc 67.0
r81 n109 n109___rc 105.0
r82 n110 n110___rc 85.0
r83 n113 n113___rc 103.0
r84 n114 n114___rc 143.0
r85 n115 n115___rc 129.0
r86 n116 n116___rc 141.0
r87 n117 n117___rc 99.0
r88 n118 n118___rc 148.0
r89 n119 n119___rc 99.0
r90 n120 n120___rc 153.0
r91 n121 n121___rc 179.0
r92 n122 n122___rc 112.0
r93 n123 n123___rc 97.0
r94 n124 n124___rc 153.0
r95 n125 n125___rc 157.0
r96 n126 n126___rc 98.0
r97 n127 n127___rc 97.0
r98 n128 n128___rc 26.0
r99 n131 n131___rc 40.0
r100 n132 n132___rc 21.0
r101 n133 n133___rc 8.0
r102 n134 n134___rc 10.0
r103 n135 n135___rc 21.0
r104 n136 n136___rc 71.0
r105 n137 n137___rc 80.0
r106 n138 n138___rc 15.0
r107 n139 n139___rc 62.0
r108 n140 n140___rc 37.0
r109 n141 n141___rc 52.0
r110 n142 n142___rc 52.0
r111 n143 n143___rc 13.0
r112 n144 n144___rc 29.0
r113 n145 n145___rc 8.0
r114 n146 n146___rc 31.0
r115 n147 n147___rc 11.0
r116 n148 n148___rc 19.0
r117 n149 n149___rc 12.0
r118 n150 n150___rc 72.0
r119 n151 n151___rc 10.0
r120 n152 n152___rc 34.0
r121 n153 n153___rc 60.0
r122 n154 n154___rc 31.0
r123 n155 n155___rc 47.0
r124 n156 n156___rc 30.0
r125 n157 n157___rc 75.0
r126 n158 n158___rc 17.0
r127 n159 n159___rc 50.0
r128 n160 n160___rc 54.0
r129 n161 n161___rc 62.0
r130 n162 n162___rc 20.0
r131 n163 n163___rc 13.0
r132 n164 n164___rc 20.0
r133 n165 n165___rc 6.0
r134 n166 n166___rc 24.0
r135 n167 n167___rc 27.0
r136 n168 n168___rc 13.0
r137 n169 n169___rc 31.0
r138 n170 n170___rc 19.0
r139 n171 n171___rc 15.0
r140 n172 n172___rc 9.0
r141 n173 n173___rc 9.0
r142 n174 n174___rc 10.0
r143 n175 n175___rc 22.0
r144 n176 n176___rc 33.0
r145 n177 n177___rc 37.0
r146 n178 n178___rc 8.0
r147 n179 n179___rc 15.0
r148 n180 n180___rc 7.0
r149 n181 n181___rc 17.0
r150 n182 n182___rc 8.0
r151 n183 n183___rc 31.0
r152 n184 n184___rc 38.0
r153 n185 n185___rc 21.0
r154 n186 n186___rc 44.0
r155 n187 n187___rc 75.0
r156 n188 n188___rc 16.0
r157 n189 n189___rc 38.0
r158 n190 n190___rc 55.0
r159 n191 n191___rc 70.0
r160 n192 n192___rc 22.0
r161 n193 n193___rc 58.0
r162 n194 n194___rc 19.0
r163 n195 n195___rc 46.0
r164 n196 n196___rc 41.0
r165 n197 n197___rc 27.0
r166 n198 n198___rc 23.0
r167 n199 n199___rc 29.0
r168 n200 n200___rc 22.0
r169 n201 n201___rc 17.0
r170 n202 n202___rc 36.0
r171 n203 n203___rc 25.0
r172 n204 n204___rc 32.0
r173 n205 n205___rc 47.0
r174 n206 n206___rc 34.0
r175 n207 n207___rc 38.0
r176 n208 n208___rc 61.0
r177 n209 n209___rc 62.0
r178 n229 n229___rc 46.0
r179 n231 n231___rc 34.0
r180 n232 n232___rc 4.0
r181 n233 n233___rc 69.0
r182 n234 n234___rc 9.0
r183 n235 n235___rc 24.0
r184 n236 n236___rc 39.0
r185 n237 n237___rc 14.0
r186 n238 n238___rc 14.0
r187 n239 n239___rc 19.0
r188 n240 n240___rc 9.0
r189 n241 n241___rc 14.0
r190 n242 n242___rc 78.0
r191 n243 n243___rc 12.0
r192 n244 n244___rc 19.0
r193 n245 n245___rc 8.0
r194 n246 n246___rc 44.0
r195 n247 n247___rc 4.0
r196 n248 n248___rc 2.0
r197 n249 n249___rc 6.0
r198 n250 n250___rc 59.0
r199 n251 n251___rc 14.0
r200 n252 n252___rc 18.0
r201 n253 n253___rc 12.0
r202 n254 n254___rc 68.0
r203 n255 n255___rc 6.0
r204 n256 n256___rc 20.0
r205 n257 n257___rc 2.0
r206 n258 n258___rc 63.0
r207 n259 n259___rc 3.0
r208 n260 n260___rc 27.0
r209 n261 n261___rc 18.0
r210 n262 n262___rc 35.0
r211 n263 n263___rc 3.0
r212 n264 n264___rc 6.0
r213 n265 n265___rc 35.0
r214 n266 n266___rc 50.0
r215 n267 n267___rc 11.0
r216 n268 n268___rc 4.0
r217 n269 n269___rc 7.0
r218 n270 n270___rc 67.0
r219 n271 n271___rc 25.0
r220 n273 n273___rc 6.0
r221 n274 n274___rc 77.0
r222 n276 n276___rc 5.0
r223 n277 n277___rc 39.0
r224 n278 n278___rc 6.0
r225 n279 n279___rc 52.0
r226 n280 n280___rc 4.0
r227 n281 n281___rc 66.0
r228 n282 n282___rc 18.0
r229 n283 n283___rc 70.0
r230 n284 n284___rc 13.0
r231 n288 n288___rc 16.0
r232 n290 n290___rc 5.0
r233 n293 n293___rc 19.0
r234 n295 n295___rc 41.0
r235 n297 n297___rc 7.0
r236 n299 n299___rc 18.0
r237 n301 n301___rc 11.0
r238 n303 n303___rc 31.0
r239 n305 n305___rc 12.0
r240 n307 n307___rc 7.0
r241 n309 n309___rc 12.0
r242 n311 n311___rc 13.0
r243 n313 n313___rc 12.0
r244 n315 n315___rc 10.0
r245 n317 n317___rc 12.0
r246 n319 n319___rc 4.0
r247 n322 n322___rc 143.0
r248 n323 n323___rc 4.0
r249 n324 n324___rc 5.0
r250 n325 n325___rc 3.0
r251 n326 n326___rc 33.0
r252 n327 n327___rc 52.0
r253 n328 n328___rc 6.0
r254 n336 n336___rc 74.0
r255 n337 n337___rc 23.0
r256 n338 n338___rc 14.0
r257 n339 n339___rc 95.0
r258 n344 n344___rc 55.0
r259 n348 n348___rc 9.0
r260 n349 n349___rc 11.0
r261 n350 n350___rc 8.0
r262 n351 n351___rc 14.0
r263 n352 n352___rc 30.0
r264 n353 n353___rc 38.0
r265 n354 n354___rc 29.0
r266 n355 n355___rc 14.0
r267 n357 n357___rc 6.0
r268 n358 n358___rc 14.0
r269 n359 n359___rc 11.0
r270 n360 n360___rc 26.0
r271 n361 n361___rc 34.0
r272 n362 n362___rc 50.0
r273 n363 n363___rc 31.0
r274 n364 n364___rc 36.0
r275 n365 n365___rc 22.0
r276 n366 n366___rc 9.0
r277 n367 n367___rc 26.0
r278 n368 n368___rc 30.0
r279 n369 n369___rc 22.0
r280 n370 n370___rc 5.0
r281 n371 n371___rc 70.0
r282 n372 n372___rc 48.0
r283 n373 n373___rc 17.0
r284 n374 n374___rc 79.0
r285 n375 n375___rc 11.0
r286 n376 n376___rc 12.0
r287 n377 n377___rc 15.0
r288 n378 n378___rc 78.0
r289 n380 n380___rc 18.0
r290 n381 n381___rc 7.0
r291 n383 n383___rc 4.0
r292 n384 n384___rc 49.0
r293 n385 n385___rc 31.0
r294 n386 n386___rc 32.0
r295 n387 n387___rc 59.0
r296 n388 n388___rc 47.0
r297 n389 n389___rc 28.0
r298 n390 n390___rc 42.0
r299 n391 n391___rc 11.0
r300 n392 n392___rc 56.0
r301 n393 n393___rc 12.0
r302 n394 n394___rc 2.0
r303 n395 n395___rc 13.0
r304 n396 n396___rc 11.0
r305 n397 n397___rc 4.0
r306 n399 n399___rc 68.0
r307 n400 n400___rc 35.0
r308 n401 n401___rc 59.0
r309 n402 n402___rc 80.0
r310 n403 n403___rc 66.0
r311 n404 n404___rc 69.0
r312 n405 n405___rc 68.0
r313 n406 n406___rc 68.0
r314 n407 n407___rc 62.0
r315 n408 n408___rc 71.0
r316 n409 n409___rc 34.0
r317 n410 n410___rc 20.0
r318 n411 n411___rc 32.0
r319 n412 n412___rc 35.0
r320 n413 n413___rc 25.0
r321 n438 n438___rc 6.0
r322 n440 n440___rc 36.0
r323 n441 n441___rc 23.0
r324 n443 n443___rc 15.0
r325 n444 n444___rc 11.0
r326 n446 n446___rc 8.0
r327 n447 n447___rc 52.0
r328 n448 n448___rc 20.0
r329 n450 n450___rc 23.0
r330 n451 n451___rc 29.0
r331 n468 n468___rc 41.0
r332 n485 n485___rc 21.0
r333 n486 n486___rc 9.0
r334 n487 n487___rc 13.0
r335 n488 n488___rc 8.0
r336 n489 n489___rc 10.0
r337 n490 n490___rc 9.0
r338 n491 n491___rc 8.0
r339 n492 n492___rc 46.0
r340 n493 n493___rc 15.0
r341 n494 n494___rc 20.0
r342 n495 n495___rc 5.0
r343 n496 n496___rc 17.0
r344 n497 n497___rc 40.0
r345 n498 n498___rc 12.0
r346 n499 n499___rc 17.0
r347 n500 n500___rc 12.0
r348 n501 n501___rc 11.0
r349 n502 n502___rc 6.0
r350 n503 n503___rc 29.0
r351 n504 n504___rc 26.0
r352 n505 n505___rc 13.0
r353 n506 n506___rc 29.0
r354 n507 n507___rc 25.0
r355 n508 n508___rc 5.0
r356 n509 n509___rc 47.0
r357 n512 n512___rc 16.0
r358 n513 n513___rc 12.0
r359 n514 n514___rc 7.0
r360 n515 n515___rc 11.0
r361 n516 n516___rc 11.0
r362 n517 n517___rc 6.0
r363 n518 n518___rc 61.0
r364 n519 n519___rc 70.0
r365 n520 n520___rc 11.0
r366 n521 n521___rc 57.0
r367 n522 n522___rc 58.0
r368 n523 n523___rc 29.0
r369 n524 n524___rc 71.0
r370 n525 n525___rc 90.0
r371 n526 n526___rc 19.0
r372 n527 n527___rc 10.0
r373 n529 n529___rc 20.0
r374 n530 n530___rc 1.0
r375 n531 n531___rc 29.0
r376 n559 n559___rc 69.0
r377 n560 n560___rc 55.0
r378 n561 n561___rc 1.0
r379 n562 n562___rc 132.0
r380 n564 n564___rc 1.0
r381 n566 n566___rc 165.0
r382 n567 n567___rc 56.0
r383 n568 n568___rc 74.0
r384 n569 n569___rc 61.0
r385 n570 n570___rc 117.0
r386 n571 n571___rc 82.0
r387 n572 n572___rc 225.0
r388 n573 n573___rc 209.0
r389 n574 n574___rc 105.0
r390 n575 n575___rc 162.0
r391 n576 n576___rc 153.0
r392 n577 n577___rc 152.0
r393 n578 n578___rc 109.0
r394 n579 n579___rc 3.0
r395 n580 n580___rc 149.0
r396 n581 n581___rc 171.0
r397 n582 n582___rc 134.0
r398 n583 n583___rc 170.0
r399 n584 n584___rc 133.0
r400 n585 n585___rc 137.0
r401 n74 n74___rc 38.0
r402 n77 n77___rc 47.0
r403 n78 n78___rc 60.0
r404 n79 n79___rc 47.0
r405 n80 n80___rc 46.0
r406 n81 n81___rc 103.0
r407 n82 n82___rc 108.0
r408 n83 n83___rc 76.0
r409 n84 n84___rc 43.0
r410 n85 n85___rc 57.0
r411 n86 n86___rc 69.0
r412 n87 n87___rc 57.0
r413 n88 n88___rc 80.0
r414 n89 n89___rc 66.0
r415 n90 n90___rc 66.0
r416 n91 n91___rc 72.0
r417 n92 n92___rc 22.0
r418 n95 n95___rc 26.0
r419 n96 n96___rc 81.0
r420 n97 n97___rc 56.0
r421 n98 n98___rc 85.0
r422 n99 n99___rc 37.0
r423 pisos_0__SP1_16_N2 pisos_0__SP1_16_N2___rc 22.0
r424 pisos_0__SP1_16_N3 pisos_0__SP1_16_N3___rc 44.0
r425 pisos_0__SP1_16_N4 pisos_0__SP1_16_N4___rc 22.0
r426 pisos_0__SP1_16_ctr_1_ pisos_0__SP1_16_ctr_1____rc 14.0
r427 pisos_0__SP1_16_ctr_2_ pisos_0__SP1_16_ctr_2____rc 19.0
r428 pisos_0__SP1_16_ctr_3_ pisos_0__SP1_16_ctr_3____rc 33.0
r429 pisos_0__SP1_16_shift_reg_10_ pisos_0__SP1_16_shift_reg_10____rc 32.0
r430 pisos_0__SP1_16_shift_reg_11_ pisos_0__SP1_16_shift_reg_11____rc 1.0
r431 pisos_0__SP1_16_shift_reg_12_ pisos_0__SP1_16_shift_reg_12____rc 37.0
r432 pisos_0__SP1_16_shift_reg_13_ pisos_0__SP1_16_shift_reg_13____rc 13.0
r433 pisos_0__SP1_16_shift_reg_14_ pisos_0__SP1_16_shift_reg_14____rc 40.0
r434 pisos_0__SP1_16_shift_reg_15_ pisos_0__SP1_16_shift_reg_15____rc 13.0
r435 pisos_0__SP1_16_shift_reg_1_ pisos_0__SP1_16_shift_reg_1____rc 3.0
r436 pisos_0__SP1_16_shift_reg_2_ pisos_0__SP1_16_shift_reg_2____rc 4.0
r437 pisos_0__SP1_16_shift_reg_3_ pisos_0__SP1_16_shift_reg_3____rc 34.0
r438 pisos_0__SP1_16_shift_reg_4_ pisos_0__SP1_16_shift_reg_4____rc 28.0
r439 pisos_0__SP1_16_shift_reg_5_ pisos_0__SP1_16_shift_reg_5____rc 39.0
r440 pisos_0__SP1_16_shift_reg_6_ pisos_0__SP1_16_shift_reg_6____rc 21.0
r441 pisos_0__SP1_16_shift_reg_7_ pisos_0__SP1_16_shift_reg_7____rc 45.0
r442 pisos_0__SP1_16_shift_reg_8_ pisos_0__SP1_16_shift_reg_8____rc 41.0
r443 pisos_0__SP1_16_shift_reg_9_ pisos_0__SP1_16_shift_reg_9____rc 29.0
r444 pisos_1__SP1_16_N2 pisos_1__SP1_16_N2___rc 36.0
r445 pisos_1__SP1_16_N3 pisos_1__SP1_16_N3___rc 21.0
r446 pisos_1__SP1_16_N4 pisos_1__SP1_16_N4___rc 14.0
r447 pisos_1__SP1_16_ctr_1_ pisos_1__SP1_16_ctr_1____rc 58.0
r448 pisos_1__SP1_16_ctr_2_ pisos_1__SP1_16_ctr_2____rc 17.0
r449 pisos_1__SP1_16_ctr_3_ pisos_1__SP1_16_ctr_3____rc 8.0
r450 pisos_1__SP1_16_shift_reg_10_ pisos_1__SP1_16_shift_reg_10____rc 15.0
r451 pisos_1__SP1_16_shift_reg_11_ pisos_1__SP1_16_shift_reg_11____rc 19.0
r452 pisos_1__SP1_16_shift_reg_12_ pisos_1__SP1_16_shift_reg_12____rc 8.0
r453 pisos_1__SP1_16_shift_reg_13_ pisos_1__SP1_16_shift_reg_13____rc 20.0
r454 pisos_1__SP1_16_shift_reg_14_ pisos_1__SP1_16_shift_reg_14____rc 7.0
r455 pisos_1__SP1_16_shift_reg_15_ pisos_1__SP1_16_shift_reg_15____rc 28.0
r456 pisos_1__SP1_16_shift_reg_1_ pisos_1__SP1_16_shift_reg_1____rc 21.0
r457 pisos_1__SP1_16_shift_reg_2_ pisos_1__SP1_16_shift_reg_2____rc 8.0
r458 pisos_1__SP1_16_shift_reg_3_ pisos_1__SP1_16_shift_reg_3____rc 25.0
r459 pisos_1__SP1_16_shift_reg_4_ pisos_1__SP1_16_shift_reg_4____rc 31.0
r460 pisos_1__SP1_16_shift_reg_5_ pisos_1__SP1_16_shift_reg_5____rc 31.0
r461 pisos_1__SP1_16_shift_reg_6_ pisos_1__SP1_16_shift_reg_6____rc 18.0
r462 pisos_1__SP1_16_shift_reg_7_ pisos_1__SP1_16_shift_reg_7____rc 42.0
r463 pisos_1__SP1_16_shift_reg_8_ pisos_1__SP1_16_shift_reg_8____rc 44.0
r464 pisos_1__SP1_16_shift_reg_9_ pisos_1__SP1_16_shift_reg_9____rc 20.0
r465 pisos_2__SP1_16_N2 pisos_2__SP1_16_N2___rc 9.0
r466 pisos_2__SP1_16_N3 pisos_2__SP1_16_N3___rc 12.0
r467 pisos_2__SP1_16_N4 pisos_2__SP1_16_N4___rc 15.0
r468 pisos_2__SP1_16_ctr_1_ pisos_2__SP1_16_ctr_1____rc 27.0
r469 pisos_2__SP1_16_ctr_2_ pisos_2__SP1_16_ctr_2____rc 13.0
r470 pisos_2__SP1_16_ctr_3_ pisos_2__SP1_16_ctr_3____rc 29.0
r471 pisos_2__SP1_16_shift_reg_10_ pisos_2__SP1_16_shift_reg_10____rc 26.0
r472 pisos_2__SP1_16_shift_reg_11_ pisos_2__SP1_16_shift_reg_11____rc 37.0
r473 pisos_2__SP1_16_shift_reg_12_ pisos_2__SP1_16_shift_reg_12____rc 18.0
r474 pisos_2__SP1_16_shift_reg_13_ pisos_2__SP1_16_shift_reg_13____rc 21.0
r475 pisos_2__SP1_16_shift_reg_14_ pisos_2__SP1_16_shift_reg_14____rc 39.0
r476 pisos_2__SP1_16_shift_reg_15_ pisos_2__SP1_16_shift_reg_15____rc 34.0
r477 pisos_2__SP1_16_shift_reg_1_ pisos_2__SP1_16_shift_reg_1____rc 6.0
r478 pisos_2__SP1_16_shift_reg_2_ pisos_2__SP1_16_shift_reg_2____rc 21.0
r479 pisos_2__SP1_16_shift_reg_3_ pisos_2__SP1_16_shift_reg_3____rc 55.0
r480 pisos_2__SP1_16_shift_reg_4_ pisos_2__SP1_16_shift_reg_4____rc 24.0
r481 pisos_2__SP1_16_shift_reg_5_ pisos_2__SP1_16_shift_reg_5____rc 11.0
r482 pisos_2__SP1_16_shift_reg_6_ pisos_2__SP1_16_shift_reg_6____rc 43.0
r483 pisos_2__SP1_16_shift_reg_7_ pisos_2__SP1_16_shift_reg_7____rc 23.0
r484 pisos_2__SP1_16_shift_reg_8_ pisos_2__SP1_16_shift_reg_8____rc 8.0
r485 pisos_2__SP1_16_shift_reg_9_ pisos_2__SP1_16_shift_reg_9____rc 20.0
r486 pisos_3__SP1_16_N1 pisos_3__SP1_16_N1___rc 14.0
r487 pisos_3__SP1_16_N2 pisos_3__SP1_16_N2___rc 48.0
r488 pisos_3__SP1_16_N3 pisos_3__SP1_16_N3___rc 8.0
r489 pisos_3__SP1_16_N4 pisos_3__SP1_16_N4___rc 19.0
r490 pisos_3__SP1_16_ctr_0_ pisos_3__SP1_16_ctr_0____rc 52.0
r491 pisos_3__SP1_16_ctr_1_ pisos_3__SP1_16_ctr_1____rc 66.0
r492 pisos_3__SP1_16_ctr_2_ pisos_3__SP1_16_ctr_2____rc 8.0
r493 pisos_3__SP1_16_ctr_3_ pisos_3__SP1_16_ctr_3____rc 19.0
r494 pisos_3__SP1_16_shift_reg_10_ pisos_3__SP1_16_shift_reg_10____rc 28.0
r495 pisos_3__SP1_16_shift_reg_11_ pisos_3__SP1_16_shift_reg_11____rc 12.0
r496 pisos_3__SP1_16_shift_reg_12_ pisos_3__SP1_16_shift_reg_12____rc 19.0
r497 pisos_3__SP1_16_shift_reg_13_ pisos_3__SP1_16_shift_reg_13____rc 37.0
r498 pisos_3__SP1_16_shift_reg_14_ pisos_3__SP1_16_shift_reg_14____rc 22.0
r499 pisos_3__SP1_16_shift_reg_15_ pisos_3__SP1_16_shift_reg_15____rc 69.0
r500 pisos_3__SP1_16_shift_reg_1_ pisos_3__SP1_16_shift_reg_1____rc 13.0
r501 pisos_3__SP1_16_shift_reg_2_ pisos_3__SP1_16_shift_reg_2____rc 41.0
r502 pisos_3__SP1_16_shift_reg_3_ pisos_3__SP1_16_shift_reg_3____rc 35.0
r503 pisos_3__SP1_16_shift_reg_4_ pisos_3__SP1_16_shift_reg_4____rc 14.0
r504 pisos_3__SP1_16_shift_reg_5_ pisos_3__SP1_16_shift_reg_5____rc 11.0
r505 pisos_3__SP1_16_shift_reg_6_ pisos_3__SP1_16_shift_reg_6____rc 21.0
r506 pisos_3__SP1_16_shift_reg_7_ pisos_3__SP1_16_shift_reg_7____rc 10.0
r507 pisos_3__SP1_16_shift_reg_8_ pisos_3__SP1_16_shift_reg_8____rc 29.0
r508 pisos_3__SP1_16_shift_reg_9_ pisos_3__SP1_16_shift_reg_9____rc 14.0
*** Estimated net capacitances from Design Compiler
c1 CLK_IN___rc VSS_SIPO4_64 5.8446e-17
c2 DATA_USED_OUT___rc VSS_SIPO4_64 6.2218e-16
c3 PARALLEL_OUT[0]___rc VSS_SIPO4_64 7.35981e-16
c4 PARALLEL_OUT[10]___rc VSS_SIPO4_64 7.88264e-16
c5 PARALLEL_OUT[11]___rc VSS_SIPO4_64 4.66151e-16
c6 PARALLEL_OUT[12]___rc VSS_SIPO4_64 5.78893e-16
c7 PARALLEL_OUT[13]___rc VSS_SIPO4_64 2.56526e-16
c8 PARALLEL_OUT[14]___rc VSS_SIPO4_64 5.21425e-16
c9 PARALLEL_OUT[15]___rc VSS_SIPO4_64 6.10891e-16
c10 PARALLEL_OUT[16]___rc VSS_SIPO4_64 2.9437e-16
c11 PARALLEL_OUT[17]___rc VSS_SIPO4_64 2.45385e-16
c12 PARALLEL_OUT[18]___rc VSS_SIPO4_64 5.81573e-16
c13 PARALLEL_OUT[19]___rc VSS_SIPO4_64 8.61891e-16
c14 PARALLEL_OUT[1]___rc VSS_SIPO4_64 7.32237e-16
c15 PARALLEL_OUT[20]___rc VSS_SIPO4_64 5.54161e-16
c16 PARALLEL_OUT[21]___rc VSS_SIPO4_64 4.8824e-16
c17 PARALLEL_OUT[22]___rc VSS_SIPO4_64 3.88937e-16
c18 PARALLEL_OUT[23]___rc VSS_SIPO4_64 8.73933e-16
c19 PARALLEL_OUT[24]___rc VSS_SIPO4_64 6.5328e-16
c20 PARALLEL_OUT[25]___rc VSS_SIPO4_64 7.45063e-16
c21 PARALLEL_OUT[26]___rc VSS_SIPO4_64 7.22973e-16
c22 PARALLEL_OUT[27]___rc VSS_SIPO4_64 8.0684e-16
c23 PARALLEL_OUT[28]___rc VSS_SIPO4_64 7.22362e-16
c24 PARALLEL_OUT[29]___rc VSS_SIPO4_64 5.35587e-16
c25 PARALLEL_OUT[2]___rc VSS_SIPO4_64 8.01258e-16
c26 PARALLEL_OUT[30]___rc VSS_SIPO4_64 6.54037e-16
c27 PARALLEL_OUT[31]___rc VSS_SIPO4_64 5.16163e-16
c28 PARALLEL_OUT[32]___rc VSS_SIPO4_64 7.48711e-16
c29 PARALLEL_OUT[33]___rc VSS_SIPO4_64 5.41512e-16
c30 PARALLEL_OUT[34]___rc VSS_SIPO4_64 7.945e-16
c31 PARALLEL_OUT[35]___rc VSS_SIPO4_64 8.51142e-16
c32 PARALLEL_OUT[36]___rc VSS_SIPO4_64 6.33979e-16
c33 PARALLEL_OUT[37]___rc VSS_SIPO4_64 3.11424e-16
c34 PARALLEL_OUT[38]___rc VSS_SIPO4_64 3.07909e-16
c35 PARALLEL_OUT[39]___rc VSS_SIPO4_64 8.58417e-16
c36 PARALLEL_OUT[3]___rc VSS_SIPO4_64 8.65623e-16
c37 PARALLEL_OUT[40]___rc VSS_SIPO4_64 7.17339e-16
c38 PARALLEL_OUT[41]___rc VSS_SIPO4_64 1.096846e-15
c39 PARALLEL_OUT[42]___rc VSS_SIPO4_64 4.84832e-16
c40 PARALLEL_OUT[43]___rc VSS_SIPO4_64 6.03656e-16
c41 PARALLEL_OUT[44]___rc VSS_SIPO4_64 2.8229e-16
c42 PARALLEL_OUT[45]___rc VSS_SIPO4_64 9.70859e-16
c43 PARALLEL_OUT[46]___rc VSS_SIPO4_64 5.64793e-16
c44 PARALLEL_OUT[47]___rc VSS_SIPO4_64 7.83527e-16
c45 PARALLEL_OUT[48]___rc VSS_SIPO4_64 7.81068e-16
c46 PARALLEL_OUT[49]___rc VSS_SIPO4_64 1.198938e-15
c47 PARALLEL_OUT[4]___rc VSS_SIPO4_64 5.79554e-16
c48 PARALLEL_OUT[50]___rc VSS_SIPO4_64 5.97743e-16
c49 PARALLEL_OUT[51]___rc VSS_SIPO4_64 1.101219e-15
c50 PARALLEL_OUT[52]___rc VSS_SIPO4_64 1.074058e-15
c51 PARALLEL_OUT[53]___rc VSS_SIPO4_64 8.96537e-16
c52 PARALLEL_OUT[54]___rc VSS_SIPO4_64 5.01828e-16
c53 PARALLEL_OUT[55]___rc VSS_SIPO4_64 5.8145e-16
c54 PARALLEL_OUT[56]___rc VSS_SIPO4_64 5.87788e-16
c55 PARALLEL_OUT[57]___rc VSS_SIPO4_64 1.007023e-15
c56 PARALLEL_OUT[58]___rc VSS_SIPO4_64 4.83109e-16
c57 PARALLEL_OUT[59]___rc VSS_SIPO4_64 6.44996e-16
c58 PARALLEL_OUT[5]___rc VSS_SIPO4_64 3.32345e-16
c59 PARALLEL_OUT[60]___rc VSS_SIPO4_64 6.94107e-16
c60 PARALLEL_OUT[61]___rc VSS_SIPO4_64 1.061507e-15
c61 PARALLEL_OUT[62]___rc VSS_SIPO4_64 1.262365e-15
c62 PARALLEL_OUT[63]___rc VSS_SIPO4_64 5.09209e-16
c63 PARALLEL_OUT[6]___rc VSS_SIPO4_64 8.83655e-16
c64 PARALLEL_OUT[7]___rc VSS_SIPO4_64 6.48182e-16
c65 PARALLEL_OUT[8]___rc VSS_SIPO4_64 6.02859e-16
c66 PARALLEL_OUT[9]___rc VSS_SIPO4_64 4.35883e-16
c67 RESET_IN___rc VSS_SIPO4_64 2.717523e-15
c68 SERIAL_IN[0]___rc VSS_SIPO4_64 1.61889e-16
c69 SERIAL_IN[1]___rc VSS_SIPO4_64 1.33047e-16
c70 SERIAL_IN[2]___rc VSS_SIPO4_64 8.5077e-17
c71 SERIAL_IN[3]___rc VSS_SIPO4_64 4.79992e-16
c72 n100___rc VSS_SIPO4_64 1.04959e-15
c73 n101___rc VSS_SIPO4_64 6.09459e-16
c74 n102___rc VSS_SIPO4_64 3.41759e-16
c75 n103___rc VSS_SIPO4_64 3.98154e-16
c76 n104___rc VSS_SIPO4_64 3.45106e-16
c77 n105___rc VSS_SIPO4_64 1.82308e-16
c78 n106___rc VSS_SIPO4_64 8.97785e-16
c79 n107___rc VSS_SIPO4_64 4.87426e-16
c80 n108___rc VSS_SIPO4_64 8.46278e-16
c81 n109___rc VSS_SIPO4_64 1.119166e-15
c82 n110___rc VSS_SIPO4_64 9.34144e-16
c83 n113___rc VSS_SIPO4_64 1.10796e-15
c84 n114___rc VSS_SIPO4_64 1.647751e-15
c85 n115___rc VSS_SIPO4_64 1.374149e-15
c86 n116___rc VSS_SIPO4_64 1.671365e-15
c87 n117___rc VSS_SIPO4_64 1.058084e-15
c88 n118___rc VSS_SIPO4_64 1.749924e-15
c89 n119___rc VSS_SIPO4_64 1.05985e-15
c90 n120___rc VSS_SIPO4_64 1.642818e-15
c91 n121___rc VSS_SIPO4_64 2.17033e-15
c92 n122___rc VSS_SIPO4_64 1.189232e-15
c93 n123___rc VSS_SIPO4_64 1.037336e-15
c94 n124___rc VSS_SIPO4_64 1.769215e-15
c95 n125___rc VSS_SIPO4_64 1.804837e-15
c96 n126___rc VSS_SIPO4_64 1.139841e-15
c97 n127___rc VSS_SIPO4_64 1.08114e-15
c98 n128___rc VSS_SIPO4_64 3.8088e-16
c99 n131___rc VSS_SIPO4_64 4.34709e-16
c100 n132___rc VSS_SIPO4_64 2.27265e-16
c101 n133___rc VSS_SIPO4_64 1.30009e-16
c102 n134___rc VSS_SIPO4_64 1.18642e-16
c103 n135___rc VSS_SIPO4_64 2.41289e-16
c104 n136___rc VSS_SIPO4_64 7.64021e-16
c105 n137___rc VSS_SIPO4_64 8.58222e-16
c106 n138___rc VSS_SIPO4_64 2.093e-16
c107 n139___rc VSS_SIPO4_64 8.094e-16
c108 n140___rc VSS_SIPO4_64 5.02977e-16
c109 n141___rc VSS_SIPO4_64 6.46623e-16
c110 n142___rc VSS_SIPO4_64 6.34814e-16
c111 n143___rc VSS_SIPO4_64 1.68064e-16
c112 n144___rc VSS_SIPO4_64 3.24307e-16
c113 n145___rc VSS_SIPO4_64 1.236e-16
c114 n146___rc VSS_SIPO4_64 4.95711e-16
c115 n147___rc VSS_SIPO4_64 1.21822e-16
c116 n148___rc VSS_SIPO4_64 2.08355e-16
c117 n149___rc VSS_SIPO4_64 1.7144e-16
c118 n150___rc VSS_SIPO4_64 9.08935e-16
c119 n151___rc VSS_SIPO4_64 1.35058e-16
c120 n152___rc VSS_SIPO4_64 4.02319e-16
c121 n153___rc VSS_SIPO4_64 8.19301e-16
c122 n154___rc VSS_SIPO4_64 4.36427e-16
c123 n155___rc VSS_SIPO4_64 6.99802e-16
c124 n156___rc VSS_SIPO4_64 4.82923e-16
c125 n157___rc VSS_SIPO4_64 8.50012e-16
c126 n158___rc VSS_SIPO4_64 2.80592e-16
c127 n159___rc VSS_SIPO4_64 5.39126e-16
c128 n160___rc VSS_SIPO4_64 5.88215e-16
c129 n161___rc VSS_SIPO4_64 6.98086e-16
c130 n162___rc VSS_SIPO4_64 2.85028e-16
c131 n163___rc VSS_SIPO4_64 1.5856e-16
c132 n164___rc VSS_SIPO4_64 3.07074e-16
c133 n165___rc VSS_SIPO4_64 9.1898e-17
c134 n166___rc VSS_SIPO4_64 3.45264e-16
c135 n167___rc VSS_SIPO4_64 4.21603e-16
c136 n168___rc VSS_SIPO4_64 2.1839e-16
c137 n169___rc VSS_SIPO4_64 4.85587e-16
c138 n170___rc VSS_SIPO4_64 2.76103e-16
c139 n171___rc VSS_SIPO4_64 1.80838e-16
c140 n172___rc VSS_SIPO4_64 1.03387e-16
c141 n173___rc VSS_SIPO4_64 1.22246e-16
c142 n174___rc VSS_SIPO4_64 1.38022e-16
c143 n175___rc VSS_SIPO4_64 2.51604e-16
c144 n176___rc VSS_SIPO4_64 3.96862e-16
c145 n177___rc VSS_SIPO4_64 4.70683e-16
c146 n178___rc VSS_SIPO4_64 9.6342e-17
c147 n179___rc VSS_SIPO4_64 2.33439e-16
c148 n180___rc VSS_SIPO4_64 8.7146e-17
c149 n181___rc VSS_SIPO4_64 2.12062e-16
c150 n182___rc VSS_SIPO4_64 1.12669e-16
c151 n183___rc VSS_SIPO4_64 5.07096e-16
c152 n184___rc VSS_SIPO4_64 4.47821e-16
c153 n185___rc VSS_SIPO4_64 2.41777e-16
c154 n186___rc VSS_SIPO4_64 4.79214e-16
c155 n187___rc VSS_SIPO4_64 8.06694e-16
c156 n188___rc VSS_SIPO4_64 2.00669e-16
c157 n189___rc VSS_SIPO4_64 4.05918e-16
c158 n190___rc VSS_SIPO4_64 6.35675e-16
c159 n191___rc VSS_SIPO4_64 7.83764e-16
c160 n192___rc VSS_SIPO4_64 2.6731e-16
c161 n193___rc VSS_SIPO4_64 6.24169e-16
c162 n194___rc VSS_SIPO4_64 3.16294e-16
c163 n195___rc VSS_SIPO4_64 6.4877e-16
c164 n196___rc VSS_SIPO4_64 5.89333e-16
c165 n197___rc VSS_SIPO4_64 4.03003e-16
c166 n198___rc VSS_SIPO4_64 3.668e-16
c167 n199___rc VSS_SIPO4_64 4.41252e-16
c168 n200___rc VSS_SIPO4_64 3.1048e-16
c169 n201___rc VSS_SIPO4_64 2.83079e-16
c170 n202___rc VSS_SIPO4_64 5.79592e-16
c171 n203___rc VSS_SIPO4_64 3.93964e-16
c172 n204___rc VSS_SIPO4_64 5.10664e-16
c173 n205___rc VSS_SIPO4_64 5.52238e-16
c174 n206___rc VSS_SIPO4_64 3.94473e-16
c175 n207___rc VSS_SIPO4_64 5.08157e-16
c176 n208___rc VSS_SIPO4_64 7.54012e-16
c177 n209___rc VSS_SIPO4_64 7.42064e-16
c178 n229___rc VSS_SIPO4_64 9.35051e-16
c179 n231___rc VSS_SIPO4_64 5.29243e-16
c180 n232___rc VSS_SIPO4_64 6.079e-17
c181 n233___rc VSS_SIPO4_64 9.44007e-16
c182 n234___rc VSS_SIPO4_64 1.29037e-16
c183 n235___rc VSS_SIPO4_64 2.72857e-16
c184 n236___rc VSS_SIPO4_64 6.08626e-16
c185 n237___rc VSS_SIPO4_64 2.10724e-16
c186 n238___rc VSS_SIPO4_64 1.92357e-16
c187 n239___rc VSS_SIPO4_64 2.33556e-16
c188 n240___rc VSS_SIPO4_64 9.8756e-17
c189 n241___rc VSS_SIPO4_64 1.49054e-16
c190 n242___rc VSS_SIPO4_64 1.244463e-15
c191 n243___rc VSS_SIPO4_64 1.24455e-16
c192 n244___rc VSS_SIPO4_64 2.14647e-16
c193 n245___rc VSS_SIPO4_64 9.1557e-17
c194 n246___rc VSS_SIPO4_64 6.98358e-16
c195 n247___rc VSS_SIPO4_64 4.9858e-17
c196 n248___rc VSS_SIPO4_64 2.5985e-17
c197 n249___rc VSS_SIPO4_64 7.2572e-17
c198 n250___rc VSS_SIPO4_64 9.43358e-16
c199 n251___rc VSS_SIPO4_64 2.10033e-16
c200 n252___rc VSS_SIPO4_64 1.9957e-16
c201 n253___rc VSS_SIPO4_64 1.57709e-16
c202 n254___rc VSS_SIPO4_64 1.053815e-15
c203 n255___rc VSS_SIPO4_64 9.304e-17
c204 n256___rc VSS_SIPO4_64 2.49801e-16
c205 n257___rc VSS_SIPO4_64 3.4178e-17
c206 n258___rc VSS_SIPO4_64 1.024603e-15
c207 n259___rc VSS_SIPO4_64 5.09e-17
c208 n260___rc VSS_SIPO4_64 4.26248e-16
c209 n261___rc VSS_SIPO4_64 2.81376e-16
c210 n262___rc VSS_SIPO4_64 5.15912e-16
c211 n263___rc VSS_SIPO4_64 4.0305e-17
c212 n264___rc VSS_SIPO4_64 8.0526e-17
c213 n265___rc VSS_SIPO4_64 3.79958e-16
c214 n266___rc VSS_SIPO4_64 8.0488e-16
c215 n267___rc VSS_SIPO4_64 1.85967e-16
c216 n268___rc VSS_SIPO4_64 4.0877e-17
c217 n269___rc VSS_SIPO4_64 1.06054e-16
c218 n270___rc VSS_SIPO4_64 1.066408e-15
c219 n271___rc VSS_SIPO4_64 2.95322e-16
c220 n273___rc VSS_SIPO4_64 6.4036e-17
c221 n274___rc VSS_SIPO4_64 1.112325e-15
c222 n276___rc VSS_SIPO4_64 7.5462e-17
c223 n277___rc VSS_SIPO4_64 6.16007e-16
c224 n278___rc VSS_SIPO4_64 8.2913e-17
c225 n279___rc VSS_SIPO4_64 7.5217e-16
c226 n280___rc VSS_SIPO4_64 5.5107e-17
c227 n281___rc VSS_SIPO4_64 9.1536e-16
c228 n282___rc VSS_SIPO4_64 1.88789e-16
c229 n283___rc VSS_SIPO4_64 1.076561e-15
c230 n284___rc VSS_SIPO4_64 1.44727e-16
c231 n288___rc VSS_SIPO4_64 1.84079e-16
c232 n290___rc VSS_SIPO4_64 6.5904e-17
c233 n293___rc VSS_SIPO4_64 2.38579e-16
c234 n295___rc VSS_SIPO4_64 4.70793e-16
c235 n297___rc VSS_SIPO4_64 8.1258e-17
c236 n299___rc VSS_SIPO4_64 2.05934e-16
c237 n301___rc VSS_SIPO4_64 1.12932e-16
c238 n303___rc VSS_SIPO4_64 4.12665e-16
c239 n305___rc VSS_SIPO4_64 1.32698e-16
c240 n307___rc VSS_SIPO4_64 9.5764e-17
c241 n309___rc VSS_SIPO4_64 1.35008e-16
c242 n311___rc VSS_SIPO4_64 1.39183e-16
c243 n313___rc VSS_SIPO4_64 1.69692e-16
c244 n315___rc VSS_SIPO4_64 1.42871e-16
c245 n317___rc VSS_SIPO4_64 1.59403e-16
c246 n319___rc VSS_SIPO4_64 5.0882e-17
c247 n322___rc VSS_SIPO4_64 3.223741e-15
c248 n323___rc VSS_SIPO4_64 4.7131e-17
c249 n324___rc VSS_SIPO4_64 8.1534e-17
c250 n325___rc VSS_SIPO4_64 4.4976e-17
c251 n326___rc VSS_SIPO4_64 3.87163e-16
c252 n327___rc VSS_SIPO4_64 6.22072e-16
c253 n328___rc VSS_SIPO4_64 7.668e-17
c254 n336___rc VSS_SIPO4_64 1.022991e-15
c255 n337___rc VSS_SIPO4_64 2.97438e-16
c256 n338___rc VSS_SIPO4_64 2.213e-16
c257 n339___rc VSS_SIPO4_64 1.899147e-15
c258 n344___rc VSS_SIPO4_64 5.94044e-16
c259 n348___rc VSS_SIPO4_64 1.01129e-16
c260 n349___rc VSS_SIPO4_64 1.3659e-16
c261 n350___rc VSS_SIPO4_64 1.16062e-16
c262 n351___rc VSS_SIPO4_64 1.64587e-16
c263 n352___rc VSS_SIPO4_64 4.56009e-16
c264 n353___rc VSS_SIPO4_64 5.45275e-16
c265 n354___rc VSS_SIPO4_64 3.77471e-16
c266 n355___rc VSS_SIPO4_64 1.66523e-16
c267 n357___rc VSS_SIPO4_64 6.405e-17
c268 n358___rc VSS_SIPO4_64 2.17868e-16
c269 n359___rc VSS_SIPO4_64 1.27207e-16
c270 n360___rc VSS_SIPO4_64 4.02535e-16
c271 n361___rc VSS_SIPO4_64 3.86621e-16
c272 n362___rc VSS_SIPO4_64 6.68438e-16
c273 n363___rc VSS_SIPO4_64 3.48979e-16
c274 n364___rc VSS_SIPO4_64 5.19728e-16
c275 n365___rc VSS_SIPO4_64 3.47533e-16
c276 n366___rc VSS_SIPO4_64 9.7424e-17
c277 n367___rc VSS_SIPO4_64 3.85421e-16
c278 n368___rc VSS_SIPO4_64 3.56308e-16
c279 n369___rc VSS_SIPO4_64 2.73701e-16
c280 n370___rc VSS_SIPO4_64 7.5364e-17
c281 n371___rc VSS_SIPO4_64 8.38462e-16
c282 n372___rc VSS_SIPO4_64 5.44354e-16
c283 n373___rc VSS_SIPO4_64 2.44813e-16
c284 n374___rc VSS_SIPO4_64 9.17464e-16
c285 n375___rc VSS_SIPO4_64 1.61907e-16
c286 n376___rc VSS_SIPO4_64 1.64021e-16
c287 n377___rc VSS_SIPO4_64 1.70566e-16
c288 n378___rc VSS_SIPO4_64 1.023044e-15
c289 n380___rc VSS_SIPO4_64 2.04464e-16
c290 n381___rc VSS_SIPO4_64 1.14337e-16
c291 n383___rc VSS_SIPO4_64 6.2875e-17
c292 n384___rc VSS_SIPO4_64 5.17809e-16
c293 n385___rc VSS_SIPO4_64 3.35569e-16
c294 n386___rc VSS_SIPO4_64 3.71643e-16
c295 n387___rc VSS_SIPO4_64 6.39049e-16
c296 n388___rc VSS_SIPO4_64 5.07992e-16
c297 n389___rc VSS_SIPO4_64 3.08995e-16
c298 n390___rc VSS_SIPO4_64 4.83829e-16
c299 n391___rc VSS_SIPO4_64 1.51079e-16
c300 n392___rc VSS_SIPO4_64 7.10201e-16
c301 n393___rc VSS_SIPO4_64 1.32215e-16
c302 n394___rc VSS_SIPO4_64 2.7964e-17
c303 n395___rc VSS_SIPO4_64 1.93207e-16
c304 n396___rc VSS_SIPO4_64 1.36924e-16
c305 n397___rc VSS_SIPO4_64 5.0116e-17
c306 n399___rc VSS_SIPO4_64 8.91555e-16
c307 n400___rc VSS_SIPO4_64 5.62557e-16
c308 n401___rc VSS_SIPO4_64 7.60109e-16
c309 n402___rc VSS_SIPO4_64 1.132932e-15
c310 n403___rc VSS_SIPO4_64 9.51627e-16
c311 n404___rc VSS_SIPO4_64 9.85622e-16
c312 n405___rc VSS_SIPO4_64 9.23819e-16
c313 n406___rc VSS_SIPO4_64 9.62395e-16
c314 n407___rc VSS_SIPO4_64 9.72352e-16
c315 n408___rc VSS_SIPO4_64 1.018869e-15
c316 n409___rc VSS_SIPO4_64 5.19363e-16
c317 n410___rc VSS_SIPO4_64 3.28292e-16
c318 n411___rc VSS_SIPO4_64 4.69954e-16
c319 n412___rc VSS_SIPO4_64 5.3356e-16
c320 n413___rc VSS_SIPO4_64 3.79557e-16
c321 n438___rc VSS_SIPO4_64 9.5798e-17
c322 n440___rc VSS_SIPO4_64 4.45999e-16
c323 n441___rc VSS_SIPO4_64 2.65891e-16
c324 n443___rc VSS_SIPO4_64 1.68166e-16
c325 n444___rc VSS_SIPO4_64 1.21426e-16
c326 n446___rc VSS_SIPO4_64 1.04231e-16
c327 n447___rc VSS_SIPO4_64 1.041113e-15
c328 n448___rc VSS_SIPO4_64 3.25983e-16
c329 n450___rc VSS_SIPO4_64 3.27137e-16
c330 n451___rc VSS_SIPO4_64 4.78492e-16
c331 n468___rc VSS_SIPO4_64 5.34241e-16
c332 n485___rc VSS_SIPO4_64 2.95355e-16
c333 n486___rc VSS_SIPO4_64 1.15331e-16
c334 n487___rc VSS_SIPO4_64 1.67946e-16
c335 n488___rc VSS_SIPO4_64 1.17772e-16
c336 n489___rc VSS_SIPO4_64 1.17321e-16
c337 n490___rc VSS_SIPO4_64 1.39224e-16
c338 n491___rc VSS_SIPO4_64 8.7703e-17
c339 n492___rc VSS_SIPO4_64 7.71372e-16
c340 n493___rc VSS_SIPO4_64 1.96021e-16
c341 n494___rc VSS_SIPO4_64 3.04936e-16
c342 n495___rc VSS_SIPO4_64 5.7665e-17
c343 n496___rc VSS_SIPO4_64 2.49257e-16
c344 n497___rc VSS_SIPO4_64 5.62259e-16
c345 n498___rc VSS_SIPO4_64 1.36435e-16
c346 n499___rc VSS_SIPO4_64 1.78083e-16
c347 n500___rc VSS_SIPO4_64 1.36396e-16
c348 n501___rc VSS_SIPO4_64 1.23851e-16
c349 n502___rc VSS_SIPO4_64 8.498e-17
c350 n503___rc VSS_SIPO4_64 3.75073e-16
c351 n504___rc VSS_SIPO4_64 3.04492e-16
c352 n505___rc VSS_SIPO4_64 1.76478e-16
c353 n506___rc VSS_SIPO4_64 3.54915e-16
c354 n507___rc VSS_SIPO4_64 2.68536e-16
c355 n508___rc VSS_SIPO4_64 5.053e-17
c356 n509___rc VSS_SIPO4_64 5.41802e-16
c357 n512___rc VSS_SIPO4_64 2.42522e-16
c358 n513___rc VSS_SIPO4_64 1.54592e-16
c359 n514___rc VSS_SIPO4_64 7.8891e-17
c360 n515___rc VSS_SIPO4_64 1.6277e-16
c361 n516___rc VSS_SIPO4_64 1.21685e-16
c362 n517___rc VSS_SIPO4_64 8.7167e-17
c363 n518___rc VSS_SIPO4_64 7.97732e-16
c364 n519___rc VSS_SIPO4_64 8.78251e-16
c365 n520___rc VSS_SIPO4_64 1.24472e-16
c366 n521___rc VSS_SIPO4_64 7.1677e-16
c367 n522___rc VSS_SIPO4_64 7.16665e-16
c368 n523___rc VSS_SIPO4_64 3.71109e-16
c369 n524___rc VSS_SIPO4_64 9.35541e-16
c370 n525___rc VSS_SIPO4_64 1.160197e-15
c371 n526___rc VSS_SIPO4_64 2.18341e-16
c372 n527___rc VSS_SIPO4_64 1.12856e-16
c373 n529___rc VSS_SIPO4_64 2.13387e-16
c374 n530___rc VSS_SIPO4_64 1.9592e-17
c375 n531___rc VSS_SIPO4_64 3.19829e-16
c376 n559___rc VSS_SIPO4_64 8.14779e-16
c377 n560___rc VSS_SIPO4_64 5.95204e-16
c378 n561___rc VSS_SIPO4_64 2.1752e-17
c379 n562___rc VSS_SIPO4_64 4.267774e-15
c380 n564___rc VSS_SIPO4_64 1.3395e-17
c381 n566___rc VSS_SIPO4_64 2.523683e-15
c382 n567___rc VSS_SIPO4_64 9.0741e-16
c383 n568___rc VSS_SIPO4_64 1.136945e-15
c384 n569___rc VSS_SIPO4_64 1.094328e-15
c385 n570___rc VSS_SIPO4_64 2.53702e-15
c386 n571___rc VSS_SIPO4_64 1.74586e-15
c387 n572___rc VSS_SIPO4_64 5.818879e-15
c388 n573___rc VSS_SIPO4_64 4.076001e-15
c389 n574___rc VSS_SIPO4_64 2.161735e-15
c390 n575___rc VSS_SIPO4_64 3.676153e-15
c391 n576___rc VSS_SIPO4_64 3.428797e-15
c392 n577___rc VSS_SIPO4_64 3.420821e-15
c393 n578___rc VSS_SIPO4_64 3.200933e-15
c394 n579___rc VSS_SIPO4_64 5.2139e-17
c395 n580___rc VSS_SIPO4_64 4.555497e-15
c396 n581___rc VSS_SIPO4_64 2.325092e-15
c397 n582___rc VSS_SIPO4_64 3.82873e-15
c398 n583___rc VSS_SIPO4_64 5.429626e-15
c399 n584___rc VSS_SIPO4_64 4.402341e-15
c400 n585___rc VSS_SIPO4_64 4.534929e-15
c401 n74___rc VSS_SIPO4_64 5.66917e-16
c402 n77___rc VSS_SIPO4_64 6.22785e-16
c403 n78___rc VSS_SIPO4_64 7.77761e-16
c404 n79___rc VSS_SIPO4_64 5.51525e-16
c405 n80___rc VSS_SIPO4_64 5.74942e-16
c406 n81___rc VSS_SIPO4_64 1.201016e-15
c407 n82___rc VSS_SIPO4_64 1.277957e-15
c408 n83___rc VSS_SIPO4_64 9.03825e-16
c409 n84___rc VSS_SIPO4_64 5.25536e-16
c410 n85___rc VSS_SIPO4_64 7.52965e-16
c411 n86___rc VSS_SIPO4_64 9.13222e-16
c412 n87___rc VSS_SIPO4_64 7.75385e-16
c413 n88___rc VSS_SIPO4_64 1.006658e-15
c414 n89___rc VSS_SIPO4_64 8.58273e-16
c415 n90___rc VSS_SIPO4_64 7.79379e-16
c416 n91___rc VSS_SIPO4_64 9.31272e-16
c417 n92___rc VSS_SIPO4_64 2.34987e-16
c418 n95___rc VSS_SIPO4_64 2.81997e-16
c419 n96___rc VSS_SIPO4_64 8.76241e-16
c420 n97___rc VSS_SIPO4_64 6.15762e-16
c421 n98___rc VSS_SIPO4_64 9.29064e-16
c422 n99___rc VSS_SIPO4_64 4.21834e-16
c423 pisos_0__SP1_16_N2___rc VSS_SIPO4_64 2.42525e-16
c424 pisos_0__SP1_16_N3___rc VSS_SIPO4_64 4.81129e-16
c425 pisos_0__SP1_16_N4___rc VSS_SIPO4_64 2.38545e-16
c426 pisos_0__SP1_16_ctr_1____rc VSS_SIPO4_64 2.03271e-16
c427 pisos_0__SP1_16_ctr_2____rc VSS_SIPO4_64 2.46951e-16
c428 pisos_0__SP1_16_ctr_3____rc VSS_SIPO4_64 3.70732e-16
c429 pisos_0__SP1_16_shift_reg_10____rc VSS_SIPO4_64 4.01185e-16
c430 pisos_0__SP1_16_shift_reg_11____rc VSS_SIPO4_64 1.5242e-17
c431 pisos_0__SP1_16_shift_reg_12____rc VSS_SIPO4_64 4.27333e-16
c432 pisos_0__SP1_16_shift_reg_13____rc VSS_SIPO4_64 1.65193e-16
c433 pisos_0__SP1_16_shift_reg_14____rc VSS_SIPO4_64 4.63408e-16
c434 pisos_0__SP1_16_shift_reg_15____rc VSS_SIPO4_64 2.06202e-16
c435 pisos_0__SP1_16_shift_reg_1____rc VSS_SIPO4_64 3.0563e-17
c436 pisos_0__SP1_16_shift_reg_2____rc VSS_SIPO4_64 4.7516e-17
c437 pisos_0__SP1_16_shift_reg_3____rc VSS_SIPO4_64 4.63777e-16
c438 pisos_0__SP1_16_shift_reg_4____rc VSS_SIPO4_64 3.60557e-16
c439 pisos_0__SP1_16_shift_reg_5____rc VSS_SIPO4_64 4.35566e-16
c440 pisos_0__SP1_16_shift_reg_6____rc VSS_SIPO4_64 2.49102e-16
c441 pisos_0__SP1_16_shift_reg_7____rc VSS_SIPO4_64 5.51528e-16
c442 pisos_0__SP1_16_shift_reg_8____rc VSS_SIPO4_64 4.7661e-16
c443 pisos_0__SP1_16_shift_reg_9____rc VSS_SIPO4_64 3.75106e-16
c444 pisos_1__SP1_16_N2___rc VSS_SIPO4_64 3.94364e-16
c445 pisos_1__SP1_16_N3___rc VSS_SIPO4_64 2.53563e-16
c446 pisos_1__SP1_16_N4___rc VSS_SIPO4_64 2.11255e-16
c447 pisos_1__SP1_16_ctr_1____rc VSS_SIPO4_64 7.2114e-16
c448 pisos_1__SP1_16_ctr_2____rc VSS_SIPO4_64 2.56223e-16
c449 pisos_1__SP1_16_ctr_3____rc VSS_SIPO4_64 1.13207e-16
c450 pisos_1__SP1_16_shift_reg_10____rc VSS_SIPO4_64 1.96748e-16
c451 pisos_1__SP1_16_shift_reg_11____rc VSS_SIPO4_64 2.28727e-16
c452 pisos_1__SP1_16_shift_reg_12____rc VSS_SIPO4_64 1.14047e-16
c453 pisos_1__SP1_16_shift_reg_13____rc VSS_SIPO4_64 2.45261e-16
c454 pisos_1__SP1_16_shift_reg_14____rc VSS_SIPO4_64 9.1433e-17
c455 pisos_1__SP1_16_shift_reg_15____rc VSS_SIPO4_64 3.65513e-16
c456 pisos_1__SP1_16_shift_reg_1____rc VSS_SIPO4_64 2.54177e-16
c457 pisos_1__SP1_16_shift_reg_2____rc VSS_SIPO4_64 1.05654e-16
c458 pisos_1__SP1_16_shift_reg_3____rc VSS_SIPO4_64 3.30139e-16
c459 pisos_1__SP1_16_shift_reg_4____rc VSS_SIPO4_64 4.1929e-16
c460 pisos_1__SP1_16_shift_reg_5____rc VSS_SIPO4_64 3.48346e-16
c461 pisos_1__SP1_16_shift_reg_6____rc VSS_SIPO4_64 2.71996e-16
c462 pisos_1__SP1_16_shift_reg_7____rc VSS_SIPO4_64 4.87507e-16
c463 pisos_1__SP1_16_shift_reg_8____rc VSS_SIPO4_64 5.1733e-16
c464 pisos_1__SP1_16_shift_reg_9____rc VSS_SIPO4_64 2.40114e-16
c465 pisos_2__SP1_16_N2___rc VSS_SIPO4_64 1.22702e-16
c466 pisos_2__SP1_16_N3___rc VSS_SIPO4_64 1.56731e-16
c467 pisos_2__SP1_16_N4___rc VSS_SIPO4_64 1.93368e-16
c468 pisos_2__SP1_16_ctr_1____rc VSS_SIPO4_64 3.78682e-16
c469 pisos_2__SP1_16_ctr_2____rc VSS_SIPO4_64 1.6583e-16
c470 pisos_2__SP1_16_ctr_3____rc VSS_SIPO4_64 3.68805e-16
c471 pisos_2__SP1_16_shift_reg_10____rc VSS_SIPO4_64 3.33066e-16
c472 pisos_2__SP1_16_shift_reg_11____rc VSS_SIPO4_64 5.0943e-16
c473 pisos_2__SP1_16_shift_reg_12____rc VSS_SIPO4_64 2.21447e-16
c474 pisos_2__SP1_16_shift_reg_13____rc VSS_SIPO4_64 2.52809e-16
c475 pisos_2__SP1_16_shift_reg_14____rc VSS_SIPO4_64 4.3482e-16
c476 pisos_2__SP1_16_shift_reg_15____rc VSS_SIPO4_64 5.41419e-16
c477 pisos_2__SP1_16_shift_reg_1____rc VSS_SIPO4_64 8.5653e-17
c478 pisos_2__SP1_16_shift_reg_2____rc VSS_SIPO4_64 3.11345e-16
c479 pisos_2__SP1_16_shift_reg_3____rc VSS_SIPO4_64 7.04461e-16
c480 pisos_2__SP1_16_shift_reg_4____rc VSS_SIPO4_64 2.89874e-16
c481 pisos_2__SP1_16_shift_reg_5____rc VSS_SIPO4_64 1.50381e-16
c482 pisos_2__SP1_16_shift_reg_6____rc VSS_SIPO4_64 4.97116e-16
c483 pisos_2__SP1_16_shift_reg_7____rc VSS_SIPO4_64 2.85562e-16
c484 pisos_2__SP1_16_shift_reg_8____rc VSS_SIPO4_64 1.04412e-16
c485 pisos_2__SP1_16_shift_reg_9____rc VSS_SIPO4_64 2.39212e-16
c486 pisos_3__SP1_16_N1___rc VSS_SIPO4_64 1.51396e-16
c487 pisos_3__SP1_16_N2___rc VSS_SIPO4_64 7.19037e-16
c488 pisos_3__SP1_16_N3___rc VSS_SIPO4_64 1.1777e-16
c489 pisos_3__SP1_16_N4___rc VSS_SIPO4_64 2.24565e-16
c490 pisos_3__SP1_16_ctr_0____rc VSS_SIPO4_64 9.73708e-16
c491 pisos_3__SP1_16_ctr_1____rc VSS_SIPO4_64 1.062883e-15
c492 pisos_3__SP1_16_ctr_2____rc VSS_SIPO4_64 1.05246e-16
c493 pisos_3__SP1_16_ctr_3____rc VSS_SIPO4_64 2.49831e-16
c494 pisos_3__SP1_16_shift_reg_10____rc VSS_SIPO4_64 3.30784e-16
c495 pisos_3__SP1_16_shift_reg_11____rc VSS_SIPO4_64 1.55528e-16
c496 pisos_3__SP1_16_shift_reg_12____rc VSS_SIPO4_64 2.38644e-16
c497 pisos_3__SP1_16_shift_reg_13____rc VSS_SIPO4_64 4.03176e-16
c498 pisos_3__SP1_16_shift_reg_14____rc VSS_SIPO4_64 2.70391e-16
c499 pisos_3__SP1_16_shift_reg_15____rc VSS_SIPO4_64 7.33887e-16
c500 pisos_3__SP1_16_shift_reg_1____rc VSS_SIPO4_64 1.99934e-16
c501 pisos_3__SP1_16_shift_reg_2____rc VSS_SIPO4_64 4.68448e-16
c502 pisos_3__SP1_16_shift_reg_3____rc VSS_SIPO4_64 4.37282e-16
c503 pisos_3__SP1_16_shift_reg_4____rc VSS_SIPO4_64 1.78444e-16
c504 pisos_3__SP1_16_shift_reg_5____rc VSS_SIPO4_64 1.56796e-16
c505 pisos_3__SP1_16_shift_reg_6____rc VSS_SIPO4_64 2.64122e-16
c506 pisos_3__SP1_16_shift_reg_7____rc VSS_SIPO4_64 1.39816e-16
c507 pisos_3__SP1_16_shift_reg_8____rc VSS_SIPO4_64 3.76479e-16
c508 pisos_3__SP1_16_shift_reg_9____rc VSS_SIPO4_64 2.13517e-16
.ENDS
*** End

