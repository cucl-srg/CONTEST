***  Written by Yury Audzevich	
*** 
***  Comments, suggestions for improvement and criticism welcome
***  E-mail:  yury.audzevich~at~cl.cam.ac.uk
*** 
*** 
***  Copyright 2003-2013, University of Cambridge, Computer Laboratory. 
***  Copyright and related rights are licensed under the Hardware License, 
***  Version 2.0 (the "License"); you may not use this file except in 
***  compliance with the License. You may obtain a copy of the License at
***  http://www.cl.cam.ac.uk/research/srg/netos/greenict/projects/contest/. 
***  Unless required by applicable law or agreed to in writing, software, 
***  hardware and materials distributed under this License is distributed 
***  on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
***  either express or implied. See the License for the specific language
***  governing permissions and limitations under the License.
*** 
*** 

***** HSPICE simulation using standard cell designs *****

***** 45nm predictive technology model (FreePDK v1.4)  Typical conditions, 1.1V, 25C *****
.include "/usr/groups/ecad/kits/commercial45_v2010_12/n45-hspice-model-TT_1V10_25.spi"

***** Standard cells netlist *****
.include "/usr/groups/ecad/kits/commercial45_v2010_12/n45-library-netlist-noparasitics.spi"

***** OPTIONS *****
.option post
.option nomod
.option co=255
* .option brief
* .option probe
.option dcon=1
.option lis_new=1
**.option captab 

***** Simulation type, timestep and length *****
.param FROM_TS = '1ps'
.param TO_TS = '80ns'

.tran FROM_TS TO_TS

***** Measurements *****
.include "POWER_SER.spi"
.include "POWER_DES.spi"

***** Optionally probe only the signals that are required to speed up simulation *****
.probe V(pvp*) V(pvn*) V(pvdd*)
.probe V(VDD*) V(VSS*)
.probe V(clk*) V(o*)
.probe V(DATA*)
.probe V(RESET*)
.probe V(SERIAL*)
.probe V(PARALLEL*)

***** Drive inputs using stimulus in "test.dsi", configure driver widths *****
.param beta = "2"
.param dsiwmin = "wmin*10"
.param dsilmin = "lmin"
.include "tempdir.stimulus/test-stim.sp"

***** Import synthesised netlist, instantiate it and connect power *****
.include "P10110.instantiation.spi"
.include "PISO10_1.spi"
.include "SIPO1_10.spi"

********************** Main MCML power supplies ****************************************
*** For power analysis use separate power supplies for SER and DES
.param cml_vdd = '0.9v' 
.param cmos_vdd = '1.1v' 

* CMOS power supply
Vpdd_cmos pvdd_cmos 0 DC 1.1v
Vgnd_all gnda 0 0.0v

*** Ser ***
Vpdd_cmos_s pvdd_cmos_ser 0 DC 1.1v

*** Des ***
Vpdd_cmos_d pvdd_cmos_des 0 DC 1.1v

**************** Digital part *************************************
Vdd_ser_cmos  VDD_PISO20_2 0 "supply"
Vss_ser_cmos  VSS_PISO20_2 0 0.0V

Vdd_des_cmos  VDD_SIPO2_20 0 "supply"
Vss_des_cmos  VSS_SIPO2_20 0 0.0V

********************* end of supply voltages  *******************************


