***  Written by Yury Audzevich
*** 
***  Comments, suggestions for improvement and criticism welcome
***  E-mail:  yury.audzevich~at~cl.cam.ac.uk
*** 
*** 
***  Copyright 2003-2013, University of Cambridge, Computer Laboratory. 
***  Copyright and related rights are licensed under the Hardware License, 
***  Version 2.0 (the "License"); you may not use this file except in 
***  compliance with the License. You may obtain a copy of the License at
***  http://www.cl.cam.ac.uk/research/srg/netos/greenict/projects/contest/. 
***  Unless required by applicable law or agreed to in writing, software, 
***  hardware and materials distributed under this License is distributed 
***  on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
***  either express or implied. See the License for the specific language
***  governing permissions and limitations under the License.
*** 
*** 


***** HSPICE simulation using standard cell library  transistors *****
*** Midswing voltage gain ***

***** 45nm predictive technology model (FreePDK v1.4),  Typical conditions, 1.1V, 25C *****
.include "cells.spi"
.include "params.spi"

**** ================================================= ***
*** OPTIONS ***
.option post
.option nomod
.option co=255
*.option brief
.option dcon=1
.option lis_new=1
**.option captab 
.option accurate


**** ================================================= ***
*** MCML PARAMETERS ***

*** displacement on time axis 
.param PARAM_DELTA = 1m

*** limits on the rotated curve
.param Vx = 0
.param VxL = 0
.param VxH = 'PARAM_MCML_SWING'

.param Vtop = 'PARAM_VDD_VOLTAGE'
.param Vbot = 'PARAM_VDD_VOLTAGE-PARAM_MCML_SWING'

************************************
*** Standard run without optimisation
.dc Vx VxL VxH 0.1m

************************************

**** ================================================= ***
*** MCML and ideal bias supplies
Vvdd VDD 0 PARAM_VDD_VOLTAGE
Vsss VSS 0 PARAM_VSS_VOLTAGE
*
Vvrefn VREFN 0 SWEEP_N_BIAS_VOLTAGE
Vvrefp VREFP 0 SWEEP_P_BIAS_VOLTAGE

**** ================================================= ***
*** Topology - multiple MCML INV instances

Xinv1av Ip In O1p O1n VDD VSS VREFP VREFN INV
Xinv2av O1p O1n O2p O2n VDD VSS VREFP VREFN INV
Xinv3av O2p O2n O3p O3n VDD VSS VREFP VREFN INV
Xinv4av O3p O3n O4p O4n VDD VSS VREFP VREFN INV
Xinv5av O4p O4n Op On VDD VSS VREFP VREFN INV

*** Add small parasitic loads on outputs to be more realistic
C1a O1p 0 CLOAD
C2a O1n 0 CLOAD
C3a O2p 0 CLOAD
C4a O2n 0 CLOAD
C5a O3p 0 CLOAD
C6a O3n 0 CLOAD
C7a O4p 0 CLOAD
C8a O4n 0 CLOAD
C9a Op 0 CLOAD
C10a On 0 CLOAD

**** ================================================= ***
EIp Ip VSS VOL = 'Vbot + Vx' 
EIn In VSS VOL = 'Vtop - Vx'


**** ================================================= ***
*** Measurements ***
**** ================================================= ***
*** need to find delta Y based on deltaX, e.g. dVout/dVin = (dVout/dt)/(dVin/dt)
*** measure relative change in Vout with respect to dt and Vin

*** MAX SWING Value
.measure DC max_I MAX V(Ip,VSS) 
.measure DC max_O1 MAX V(O1p,VSS) 
.measure DC max_O2 MAX V(O2p,VSS)
.measure DC max_O3 MAX V(O3p,VSS) 
.measure DC max_O4 MAX V(O3p,VSS)  

*** VOLTAGE SWING Value
.measure DC delta_I MAX V(Ip,In)
.measure DC delta_O1 MAX V(O1p,O1n)
.measure DC delta_O2 MAX V(O2p,O2n)
.measure DC delta_O3 MAX V(O3p,O3n)
.measure DC delta_O4 MAX V(O4p,O4n)

*** MIDSWING Voltage Value
.measure mid_I Param='max_I - (delta_I/2)'
.measure mid_O1 Param='max_O1 - (delta_O1/2)'
.measure mid_O2 Param='max_O2 - (delta_O2/2)'
.measure mid_O3 Param='max_O3 - (delta_O3/2)'
.measure mid_O4 Param='max_O4 - (delta_O4/2)'

*** relative analysis -- measure value of O2p when O1p at a certain time point and value
*** inv 1 '0->1' transition
.MEAS DC REL_O2PM FIND PAR('V(O2p)') WHEN V(O1p)='mid_O1-PARAM_DELTA' RISE=LAST
.MEAS DC REL_O2PP FIND PAR('V(O2p)') WHEN V(O1p)='mid_O1+PARAM_DELTA' RISE=LAST
*** inv 1 '1->0' transition
.MEAS DC REL_O2MM FIND PAR('V(O2n)') WHEN V(O1n)='mid_O1-PARAM_DELTA' FALL=LAST
.MEAS DC REL_O2MP FIND PAR('V(O2n)') WHEN V(O1n)='mid_O1+PARAM_DELTA' FALL=LAST

*** inv 2 '0->1' transition
.MEAS DC REL_O3PM FIND PAR('V(O3p)') WHEN V(O2p)='mid_O2-PARAM_DELTA' RISE=LAST
.MEAS DC REL_O3PP FIND PAR('V(O3p)') WHEN V(O2p)='mid_O2+PARAM_DELTA' RISE=LAST
*** inv 2 '1->0' transition
.MEAS DC REL_O3MM FIND PAR('V(O3n)') WHEN V(O2n)='mid_O2-PARAM_DELTA' FALL=LAST
.MEAS DC REL_O3MP FIND PAR('V(O3n)') WHEN V(O2n)='mid_O2+PARAM_DELTA' FALL=LAST

*** inv 3 '0->1' transition
.MEAS DC REL_O4PM FIND PAR('V(O4p)') WHEN V(O3p)='mid_O3-PARAM_DELTA' RISE=LAST
.MEAS DC REL_O4PP FIND PAR('V(O4p)') WHEN V(O3p)='mid_O3+PARAM_DELTA' RISE=LAST
*** inv 3 '1->0' transition
.MEAS DC REL_O4MM FIND PAR('V(O4n)') WHEN V(O3n)='mid_O3-PARAM_DELTA' FALL=LAST
.MEAS DC REL_O4MP FIND PAR('V(O4n)') WHEN V(O3n)='mid_O3+PARAM_DELTA' FALL=LAST

*** inv 4 '0->1' transition
.MEAS DC REL_O5PM FIND PAR('V(Op)') WHEN V(O4p)='mid_O4-PARAM_DELTA' RISE=LAST
.MEAS DC REL_O5PP FIND PAR('V(Op)') WHEN V(O4p)='mid_O4+PARAM_DELTA' RISE=LAST
*** inv 4 '1->0' transition
.MEAS DC REL_O5MM FIND PAR('V(On)') WHEN V(O4n)='mid_O4-PARAM_DELTA' FALL=LAST
.MEAS DC REL_O5MP FIND PAR('V(On)') WHEN V(O4n)='mid_O4+PARAM_DELTA' FALL=LAST

*** Record the parameters in the .mt0 file
.meas DELIM0 param='0.0'
.meas dc result_vdd param='PARAM_VDD_VOLTAGE'
.meas dc result_vss param='PARAM_VSS_VOLTAGE'
.meas dc result_pulldown_width param='SWEEP_N_WIDTH'
.meas dc result_pulldown_length param='SWEEP_N_LENGTH'
.meas dc result_pullup_width param='SWEEP_P_WIDTH'
.meas dc result_pullup_length param='SWEEP_P_LENGTH'
.meas dc result_sink_width param='PARAM_NSOURCE_WIDTH'
.meas dc result_sink_length param='PARAM_NSOURCE_LENGTH'
.meas dc result_n_bias param='SWEEP_N_BIAS_VOLTAGE'
.meas dc result_p_bias param='SWEEP_P_BIAS_VOLTAGE'
.meas DELIM3 param='0.0'
.meas DELIM4 param='0.0'
.meas DELIM5 param='0.0'
.meas dc result_voltage_swing param='PARAM_MCML_SWING'
.meas dc MIDSW_GAINP_INV1 param='(REL_O2PP-REL_O2PM)/(2*PARAM_DELTA)'
.meas dc MIDSW_GAINN_INV1 param='(REL_O2MP-REL_O2MM)/(2*PARAM_DELTA)'
.meas dc MIDSW_GAINP_INV2 param='(REL_O3PP-REL_O3PM)/(2*PARAM_DELTA)'
.meas dc MIDSW_GAINN_INV2 param='(REL_O3MP-REL_O3MM)/(2*PARAM_DELTA)'
.meas dc MIDSW_GAINP_INV3 param='(REL_O4PP-REL_O4PM)/(2*PARAM_DELTA)'
.meas dc MIDSW_GAINN_INV3 param='(REL_O4MP-REL_O4MM)/(2*PARAM_DELTA)'
.meas dc MIDSW_GAINP_INV4 param='(REL_O5PP-REL_O5PM)/(2*PARAM_DELTA)'
.meas dc MIDSW_GAINN_INV4 param='(REL_O5MP-REL_O5MM)/(2*PARAM_DELTA)'
.meas dc MIDSWING_GAIN_AVG param = '(MIDSW_GAINP_INV1+MIDSW_GAINN_INV1+MIDSW_GAINP_INV2+MIDSW_GAINN_INV2+MIDSW_GAINP_INV3+MIDSW_GAINN_INV3+MIDSW_GAINP_INV4+MIDSW_GAINN_INV4)/8'

