***  Written by Yury Audzevich
*** 
***  Comments, suggestions for improvement and criticism welcome
***  E-mail:  yury.audzevich~at~cl.cam.ac.uk
*** 
*** 
***  Copyright 2003-2013, University of Cambridge, Computer Laboratory. 
***  Copyright and related rights are licensed under the Hardware License, 
***  Version 2.0 (the "License"); you may not use this file except in 
***  compliance with the License. You may obtain a copy of the License at
***  http://www.cl.cam.ac.uk/research/srg/netos/greenict/projects/contest/. 
***  Unless required by applicable law or agreed to in writing, software, 
***  hardware and materials distributed under this License is distributed 
***  on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
***  either express or implied. See the License for the specific language
***  governing permissions and limitations under the License.
*** 
*** 

*** 45nm predictive technology model (FreePDK v1.4),  Typical conditions, 1.1V, 25C ***

********************************************************************************
*** This file contains a collection of Design Parameters used in both: 	     ***
*** 1) optimization of single-level MCML logic 				     ***	
*** 2) post-opt. standard single-level MCML logic TRAN/DC type of analysis   *** 	
********************************************************************************

*** MAIN PARAMETERS ***

*** Optimization ON/OFF ('1'/'0')  ***
.param OPT_PARAM_ON = 0

*** simulation time
.param PARAM_TIME_S = 0.1ps
.param PARAM_TIME_E = 10ns

*** measurement time
.param PARAM_MEAS_S = 100ps
.param PARAM_MEAS_E = 10ns

*** supply voltages
.param PARAM_MCML_SWING = 0.4
*.param PARAM_MCML_SWING = optw(0.2, 0.2, 0.45, 0.01)

.param PARAM_CMOS_VDD_VOLTAGE = 1.1
.param PARAM_VDD_VOLTAGE = 0.9
.param PARAM_VSS_VOLTAGE = 0.0

*** derived parameters
.param PARAM_MCML_MID = '(PARAM_VDD_VOLTAGE + (PARAM_VDD_VOLTAGE-PARAM_MCML_SWING))/2'
.param PARAM_MCML_HALF_SWING = 'PARAM_MCML_SWING/2' 

*** parasitic capacitance
.param CLOAD = 0.05fF 

*** check for FANOUT ***
.param FANOUT_ON = 0

*** Define parameters to optimise and the ones to have fixed - the format is optw(initial, min, max, step)
*** In general HSPICE is more successful with fewer parameters to optimise when circuit has nonlinear responses to small deltas

*** Please comment/uncomment parameters that are needed for opt (2-4 parameters at a time for speed) ***
*** pull-up network
.param SWEEP_P_WIDTH = 0.25U
*.param SWEEP_P_WIDTH = optw(0.3U, 0.3U, 1.2U, 0.001U)
*
.param SWEEP_P_LENGTH = 0.055U
*.param SWEEP_P_LENGTH = optw(lmin, lmin, 0.5U, 0.005U)

*** pull-down
.param SWEEP_N_WIDTH = 0.21U
*.param SWEEP_N_WIDTH = optw(0.3U, wmin, 1.2U, 0.001U)
*
.param SWEEP_N_LENGTH = 'lmin'
*.param SWEEP_N_LENGTH = optw(lmin, lmin, 0.5U, 0.005U)

*** current sink 
.param PARAM_NSOURCE_WIDTH = 1.2U
*.param PARAM_NSOURCE_WIDTH = optw(1.0U, 1.0U, 3.0U, 0.001U)
*
.param PARAM_NSOURCE_LENGTH = 0.12U
*.param PARAM_NSOURCE_LENGTH = optw(lmin, lmin, 0.5U, 0.005U) 

*** reference voltages
.param SWEEP_N_BIAS_VOLTAGE = 0.53V
*.param SWEEP_N_BIAS_VOLTAGE = optw(0.3, 0.3, 0.735, 0.001)
*
.param SWEEP_P_BIAS_VOLTAGE = 50mV
*.param SWEEP_P_BIAS_VOLTAGE = optw(50m, 1m, 150m , 1m)

**** CMOS gate dimentions optimization ******
*.param SWEEP_CMOSP_WIDTH = optw(0.2U, 0.2U, 0.8U, 0.001U)
.param SWEEP_CMOSP_WIDTH = 0.3U

*.param SWEEP_CMOSN_WIDTH = optw(0.2U, 0.2U, 0.4U, 0.001U)
.param SWEEP_CMOSN_WIDTH = 0.21U




